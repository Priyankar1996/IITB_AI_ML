-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity concat is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity concat;
architecture concat_arch of concat is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal concat_CP_34_start: Boolean;
  signal concat_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ptr_deref_743_store_0_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_677_inst_req_1 : boolean;
  signal type_cast_627_inst_ack_1 : boolean;
  signal addr_of_900_final_reg_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_0 : boolean;
  signal ptr_deref_526_store_0_ack_1 : boolean;
  signal ptr_deref_526_store_0_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_695_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_677_inst_req_0 : boolean;
  signal type_cast_627_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_25_inst_ack_1 : boolean;
  signal type_cast_30_inst_req_0 : boolean;
  signal type_cast_30_inst_ack_0 : boolean;
  signal type_cast_30_inst_req_1 : boolean;
  signal type_cast_30_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_0 : boolean;
  signal type_cast_627_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_39_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_695_inst_ack_0 : boolean;
  signal type_cast_43_inst_req_0 : boolean;
  signal type_cast_627_inst_req_0 : boolean;
  signal type_cast_43_inst_ack_0 : boolean;
  signal type_cast_43_inst_req_1 : boolean;
  signal array_obj_ref_899_index_offset_req_1 : boolean;
  signal type_cast_43_inst_ack_1 : boolean;
  signal if_stmt_757_branch_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_ack_1 : boolean;
  signal call_stmt_768_call_ack_1 : boolean;
  signal type_cast_983_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_51_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_695_inst_req_0 : boolean;
  signal type_cast_55_inst_req_0 : boolean;
  signal type_cast_999_inst_req_1 : boolean;
  signal type_cast_55_inst_ack_0 : boolean;
  signal type_cast_55_inst_req_1 : boolean;
  signal type_cast_55_inst_ack_1 : boolean;
  signal type_cast_953_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_req_0 : boolean;
  signal addr_of_900_final_reg_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_0 : boolean;
  signal ptr_deref_743_store_0_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_64_inst_ack_1 : boolean;
  signal type_cast_645_inst_ack_1 : boolean;
  signal type_cast_983_inst_req_0 : boolean;
  signal type_cast_68_inst_req_0 : boolean;
  signal array_obj_ref_899_index_offset_ack_1 : boolean;
  signal type_cast_68_inst_ack_0 : boolean;
  signal type_cast_68_inst_req_1 : boolean;
  signal type_cast_68_inst_ack_1 : boolean;
  signal W_arrayidx252_894_delayed_6_0_905_inst_req_1 : boolean;
  signal type_cast_645_inst_req_1 : boolean;
  signal ptr_deref_743_store_0_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_76_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_713_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_713_inst_req_1 : boolean;
  signal type_cast_983_inst_ack_0 : boolean;
  signal type_cast_80_inst_req_0 : boolean;
  signal type_cast_80_inst_ack_0 : boolean;
  signal type_cast_80_inst_req_1 : boolean;
  signal type_cast_80_inst_ack_1 : boolean;
  signal W_arrayidx252_894_delayed_6_0_905_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_89_inst_ack_1 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0 : boolean;
  signal addr_of_607_final_reg_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_713_inst_ack_0 : boolean;
  signal type_cast_93_inst_req_0 : boolean;
  signal type_cast_93_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_ack_0 : boolean;
  signal type_cast_93_inst_req_1 : boolean;
  signal type_cast_999_inst_ack_1 : boolean;
  signal type_cast_93_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_731_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_731_inst_req_1 : boolean;
  signal type_cast_645_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_101_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_713_inst_req_0 : boolean;
  signal type_cast_645_inst_req_0 : boolean;
  signal addr_of_607_final_reg_req_1 : boolean;
  signal type_cast_105_inst_req_0 : boolean;
  signal type_cast_105_inst_ack_0 : boolean;
  signal type_cast_105_inst_req_1 : boolean;
  signal type_cast_105_inst_ack_1 : boolean;
  signal array_obj_ref_899_index_offset_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_0 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_114_inst_ack_1 : boolean;
  signal type_cast_953_inst_req_0 : boolean;
  signal type_cast_118_inst_req_0 : boolean;
  signal type_cast_118_inst_ack_0 : boolean;
  signal type_cast_118_inst_req_1 : boolean;
  signal type_cast_118_inst_ack_1 : boolean;
  signal type_cast_999_inst_ack_0 : boolean;
  signal type_cast_663_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_623_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_0 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_126_inst_ack_1 : boolean;
  signal W_arrayidx252_894_delayed_6_0_905_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_623_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_731_inst_ack_0 : boolean;
  signal type_cast_130_inst_req_0 : boolean;
  signal type_cast_130_inst_ack_0 : boolean;
  signal type_cast_130_inst_req_1 : boolean;
  signal type_cast_130_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_731_inst_req_0 : boolean;
  signal type_cast_663_inst_req_1 : boolean;
  signal type_cast_968_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_139_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_ack_1 : boolean;
  signal addr_of_900_final_reg_req_1 : boolean;
  signal type_cast_410_inst_req_0 : boolean;
  signal type_cast_410_inst_ack_0 : boolean;
  signal type_cast_410_inst_req_1 : boolean;
  signal type_cast_410_inst_ack_1 : boolean;
  signal type_cast_717_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_659_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_424_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_424_inst_ack_0 : boolean;
  signal type_cast_143_inst_req_0 : boolean;
  signal type_cast_143_inst_ack_0 : boolean;
  signal type_cast_143_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_623_inst_ack_0 : boolean;
  signal type_cast_143_inst_ack_1 : boolean;
  signal if_stmt_757_branch_req_0 : boolean;
  signal type_cast_968_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_623_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_151_inst_ack_1 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal type_cast_663_inst_ack_0 : boolean;
  signal type_cast_663_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_0 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_164_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_ack_1 : boolean;
  signal addr_of_607_final_reg_ack_0 : boolean;
  signal type_cast_168_inst_req_0 : boolean;
  signal type_cast_168_inst_ack_0 : boolean;
  signal type_cast_168_inst_req_1 : boolean;
  signal type_cast_168_inst_ack_1 : boolean;
  signal do_while_stmt_817_branch_req_0 : boolean;
  signal if_stmt_1654_branch_ack_1 : boolean;
  signal MUX_1253_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_0 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_176_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_1 : boolean;
  signal call_stmt_768_call_req_1 : boolean;
  signal type_cast_968_inst_req_1 : boolean;
  signal addr_of_607_final_reg_req_0 : boolean;
  signal type_cast_180_inst_req_0 : boolean;
  signal type_cast_180_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_req_1 : boolean;
  signal type_cast_180_inst_req_1 : boolean;
  signal type_cast_180_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_189_inst_ack_1 : boolean;
  signal addr_of_900_final_reg_req_0 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal type_cast_681_inst_ack_1 : boolean;
  signal type_cast_193_inst_req_0 : boolean;
  signal type_cast_193_inst_ack_0 : boolean;
  signal type_cast_193_inst_req_1 : boolean;
  signal type_cast_193_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_201_inst_ack_1 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal W_arrayidx252_894_delayed_6_0_905_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0 : boolean;
  signal type_cast_983_inst_ack_1 : boolean;
  signal type_cast_681_inst_req_1 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal type_cast_968_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_214_inst_ack_1 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_req_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal ptr_deref_526_store_0_ack_0 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_226_inst_ack_1 : boolean;
  signal type_cast_735_inst_ack_1 : boolean;
  signal call_stmt_768_call_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_641_inst_ack_1 : boolean;
  signal type_cast_230_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_1 : boolean;
  signal type_cast_230_inst_ack_0 : boolean;
  signal type_cast_230_inst_req_1 : boolean;
  signal type_cast_230_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_641_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_req_0 : boolean;
  signal type_cast_614_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_ack_0 : boolean;
  signal type_cast_953_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_239_inst_ack_1 : boolean;
  signal call_stmt_768_call_req_0 : boolean;
  signal type_cast_681_inst_ack_0 : boolean;
  signal type_cast_243_inst_req_0 : boolean;
  signal type_cast_243_inst_ack_0 : boolean;
  signal type_cast_681_inst_req_0 : boolean;
  signal type_cast_243_inst_req_1 : boolean;
  signal type_cast_243_inst_ack_1 : boolean;
  signal type_cast_735_inst_req_1 : boolean;
  signal type_cast_735_inst_ack_0 : boolean;
  signal type_cast_735_inst_req_0 : boolean;
  signal type_cast_953_inst_req_1 : boolean;
  signal ptr_deref_526_store_0_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_req_0 : boolean;
  signal if_stmt_308_branch_req_0 : boolean;
  signal if_stmt_308_branch_ack_1 : boolean;
  signal if_stmt_308_branch_ack_0 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0 : boolean;
  signal if_stmt_323_branch_req_0 : boolean;
  signal if_stmt_323_branch_ack_1 : boolean;
  signal if_stmt_323_branch_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_641_inst_ack_0 : boolean;
  signal type_cast_360_inst_req_0 : boolean;
  signal type_cast_360_inst_ack_0 : boolean;
  signal type_cast_360_inst_req_1 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal type_cast_360_inst_ack_1 : boolean;
  signal type_cast_717_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_677_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_641_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_659_inst_ack_1 : boolean;
  signal array_obj_ref_389_index_offset_req_0 : boolean;
  signal array_obj_ref_389_index_offset_ack_0 : boolean;
  signal array_obj_ref_389_index_offset_req_1 : boolean;
  signal array_obj_ref_389_index_offset_ack_1 : boolean;
  signal if_stmt_757_branch_ack_0 : boolean;
  signal ptr_deref_743_store_0_ack_1 : boolean;
  signal addr_of_390_final_reg_req_0 : boolean;
  signal addr_of_390_final_reg_ack_0 : boolean;
  signal addr_of_390_final_reg_req_1 : boolean;
  signal addr_of_390_final_reg_ack_1 : boolean;
  signal type_cast_717_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_659_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_ack_0 : boolean;
  signal if_stmt_540_branch_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_ack_1 : boolean;
  signal type_cast_397_inst_req_0 : boolean;
  signal type_cast_397_inst_ack_0 : boolean;
  signal type_cast_397_inst_req_1 : boolean;
  signal type_cast_397_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_424_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_424_inst_ack_1 : boolean;
  signal array_obj_ref_606_index_offset_ack_1 : boolean;
  signal type_cast_428_inst_req_0 : boolean;
  signal type_cast_428_inst_ack_0 : boolean;
  signal type_cast_428_inst_req_1 : boolean;
  signal type_cast_428_inst_ack_1 : boolean;
  signal type_cast_717_inst_req_0 : boolean;
  signal type_cast_1270_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_659_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_442_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_442_inst_ack_0 : boolean;
  signal if_stmt_540_branch_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_442_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_442_inst_ack_1 : boolean;
  signal ptr_deref_910_store_0_ack_0 : boolean;
  signal array_obj_ref_606_index_offset_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_677_inst_ack_1 : boolean;
  signal array_obj_ref_899_index_offset_req_0 : boolean;
  signal type_cast_446_inst_req_0 : boolean;
  signal type_cast_446_inst_ack_0 : boolean;
  signal type_cast_446_inst_req_1 : boolean;
  signal type_cast_446_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_460_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_460_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_460_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_460_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0 : boolean;
  signal type_cast_464_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_1 : boolean;
  signal type_cast_464_inst_ack_0 : boolean;
  signal type_cast_464_inst_req_1 : boolean;
  signal type_cast_464_inst_ack_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_478_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_478_inst_ack_0 : boolean;
  signal if_stmt_540_branch_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_478_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_478_inst_ack_1 : boolean;
  signal array_obj_ref_606_index_offset_ack_0 : boolean;
  signal array_obj_ref_606_index_offset_req_0 : boolean;
  signal type_cast_482_inst_req_0 : boolean;
  signal type_cast_482_inst_ack_0 : boolean;
  signal type_cast_482_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_610_inst_req_1 : boolean;
  signal type_cast_482_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_496_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_496_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_496_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_496_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_695_inst_ack_1 : boolean;
  signal type_cast_500_inst_req_0 : boolean;
  signal type_cast_500_inst_ack_0 : boolean;
  signal type_cast_500_inst_req_1 : boolean;
  signal type_cast_500_inst_ack_1 : boolean;
  signal ptr_deref_910_store_0_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_514_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_514_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_514_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_514_inst_ack_1 : boolean;
  signal type_cast_518_inst_req_0 : boolean;
  signal type_cast_518_inst_ack_0 : boolean;
  signal type_cast_518_inst_req_1 : boolean;
  signal type_cast_518_inst_ack_1 : boolean;
  signal phi_stmt_819_req_0 : boolean;
  signal type_cast_1073_inst_req_0 : boolean;
  signal phi_stmt_819_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0 : boolean;
  signal phi_stmt_819_ack_0 : boolean;
  signal type_cast_1036_inst_ack_1 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_999_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal type_cast_1073_inst_req_1 : boolean;
  signal type_cast_1324_inst_req_1 : boolean;
  signal phi_stmt_594_req_0 : boolean;
  signal type_cast_1298_inst_req_1 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_ack_1 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_req_1 : boolean;
  signal type_cast_1036_inst_req_1 : boolean;
  signal phi_stmt_824_req_0 : boolean;
  signal type_cast_1036_inst_ack_0 : boolean;
  signal type_cast_1036_inst_req_0 : boolean;
  signal phi_stmt_824_req_1 : boolean;
  signal phi_stmt_824_ack_0 : boolean;
  signal type_cast_827_inst_req_0 : boolean;
  signal type_cast_827_inst_ack_0 : boolean;
  signal type_cast_827_inst_req_1 : boolean;
  signal type_cast_827_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_ack_1 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_ack_0 : boolean;
  signal W_add_outx_x1_914_delayed_1_0_933_inst_req_0 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1 : boolean;
  signal do_while_stmt_817_branch_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1 : boolean;
  signal phi_stmt_829_req_0 : boolean;
  signal phi_stmt_829_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0 : boolean;
  signal type_cast_1242_inst_req_0 : boolean;
  signal phi_stmt_829_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1 : boolean;
  signal type_cast_1242_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal MUX_1253_inst_req_1 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1 : boolean;
  signal type_cast_1617_inst_ack_1 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal type_cast_1298_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0 : boolean;
  signal phi_stmt_834_req_0 : boolean;
  signal MUX_1331_inst_ack_1 : boolean;
  signal MUX_1305_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1 : boolean;
  signal phi_stmt_834_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_req_1 : boolean;
  signal phi_stmt_834_ack_0 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal MUX_1253_inst_ack_1 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal type_cast_837_inst_req_1 : boolean;
  signal type_cast_837_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0 : boolean;
  signal MUX_1305_inst_ack_0 : boolean;
  signal type_cast_1073_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0 : boolean;
  signal W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1 : boolean;
  signal MUX_1253_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0 : boolean;
  signal type_cast_1270_inst_req_1 : boolean;
  signal phi_stmt_839_req_0 : boolean;
  signal type_cast_1073_inst_ack_0 : boolean;
  signal MUX_1331_inst_req_1 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0 : boolean;
  signal phi_stmt_839_req_1 : boolean;
  signal phi_stmt_839_ack_0 : boolean;
  signal type_cast_1324_inst_ack_1 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0 : boolean;
  signal W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1625_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1 : boolean;
  signal W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0 : boolean;
  signal ptr_deref_910_store_0_ack_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1 : boolean;
  signal ptr_deref_910_store_0_req_1 : boolean;
  signal MUX_1305_inst_ack_1 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0 : boolean;
  signal W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1 : boolean;
  signal W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0 : boolean;
  signal W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0 : boolean;
  signal type_cast_1242_inst_req_1 : boolean;
  signal type_cast_870_inst_req_0 : boolean;
  signal type_cast_870_inst_ack_0 : boolean;
  signal type_cast_870_inst_req_1 : boolean;
  signal type_cast_870_inst_ack_1 : boolean;
  signal array_obj_ref_876_index_offset_req_0 : boolean;
  signal array_obj_ref_876_index_offset_ack_0 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal array_obj_ref_876_index_offset_req_1 : boolean;
  signal array_obj_ref_876_index_offset_ack_1 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal type_cast_1242_inst_ack_1 : boolean;
  signal addr_of_877_final_reg_req_0 : boolean;
  signal addr_of_877_final_reg_ack_0 : boolean;
  signal addr_of_877_final_reg_req_1 : boolean;
  signal addr_of_877_final_reg_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_ack_0 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1 : boolean;
  signal W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1 : boolean;
  signal if_stmt_1654_branch_req_0 : boolean;
  signal ptr_deref_885_load_0_req_0 : boolean;
  signal ptr_deref_885_load_0_ack_0 : boolean;
  signal ptr_deref_885_load_0_req_1 : boolean;
  signal ptr_deref_885_load_0_ack_1 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_req_0 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_ack_0 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_req_1 : boolean;
  signal W_add_outx_x1_883_delayed_1_0_887_inst_ack_1 : boolean;
  signal type_cast_893_inst_req_0 : boolean;
  signal type_cast_893_inst_ack_0 : boolean;
  signal type_cast_893_inst_req_1 : boolean;
  signal type_cast_893_inst_ack_1 : boolean;
  signal type_cast_600_inst_ack_1 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_0 : boolean;
  signal type_cast_1298_inst_ack_0 : boolean;
  signal type_cast_1298_inst_req_0 : boolean;
  signal MUX_1305_inst_req_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_0 : boolean;
  signal array_obj_ref_1079_index_offset_ack_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_1 : boolean;
  signal array_obj_ref_1079_index_offset_ack_1 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal type_cast_1246_inst_ack_1 : boolean;
  signal addr_of_1080_final_reg_req_0 : boolean;
  signal addr_of_1080_final_reg_ack_0 : boolean;
  signal addr_of_1080_final_reg_req_1 : boolean;
  signal addr_of_1080_final_reg_ack_1 : boolean;
  signal type_cast_1324_inst_ack_0 : boolean;
  signal MUX_1331_inst_ack_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_1 : boolean;
  signal W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_1 : boolean;
  signal if_stmt_1359_branch_req_0 : boolean;
  signal type_cast_1324_inst_req_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal type_cast_1294_inst_ack_1 : boolean;
  signal ptr_deref_1088_load_0_req_0 : boolean;
  signal type_cast_1294_inst_req_1 : boolean;
  signal ptr_deref_1088_load_0_ack_0 : boolean;
  signal ptr_deref_1088_load_0_req_1 : boolean;
  signal ptr_deref_1088_load_0_ack_1 : boolean;
  signal MUX_1331_inst_req_0 : boolean;
  signal type_cast_1294_inst_ack_0 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1 : boolean;
  signal W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1 : boolean;
  signal do_while_stmt_817_branch_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_req_0 : boolean;
  signal type_cast_1096_inst_req_0 : boolean;
  signal type_cast_1096_inst_ack_0 : boolean;
  signal type_cast_1096_inst_req_1 : boolean;
  signal type_cast_1617_inst_req_1 : boolean;
  signal type_cast_1096_inst_ack_1 : boolean;
  signal type_cast_1294_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1640_inst_ack_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal array_obj_ref_1102_index_offset_req_0 : boolean;
  signal array_obj_ref_1102_index_offset_ack_0 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal array_obj_ref_1102_index_offset_req_1 : boolean;
  signal array_obj_ref_1102_index_offset_ack_1 : boolean;
  signal type_cast_1246_inst_req_1 : boolean;
  signal addr_of_1103_final_reg_req_0 : boolean;
  signal addr_of_1103_final_reg_ack_0 : boolean;
  signal addr_of_1103_final_reg_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_req_0 : boolean;
  signal addr_of_1103_final_reg_ack_1 : boolean;
  signal W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_1 : boolean;
  signal type_cast_1607_inst_req_0 : boolean;
  signal W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_1 : boolean;
  signal MUX_1281_inst_ack_1 : boolean;
  signal MUX_1281_inst_req_1 : boolean;
  signal W_arrayidx278_1043_delayed_6_0_1108_inst_req_0 : boolean;
  signal W_arrayidx278_1043_delayed_6_0_1108_inst_ack_0 : boolean;
  signal W_arrayidx278_1043_delayed_6_0_1108_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_0 : boolean;
  signal W_arrayidx278_1043_delayed_6_0_1108_inst_ack_1 : boolean;
  signal if_stmt_1654_branch_ack_0 : boolean;
  signal type_cast_1246_inst_ack_0 : boolean;
  signal type_cast_1246_inst_req_0 : boolean;
  signal MUX_1281_inst_ack_0 : boolean;
  signal MUX_1281_inst_req_0 : boolean;
  signal type_cast_1274_inst_ack_1 : boolean;
  signal type_cast_1274_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_req_1 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal ptr_deref_1113_store_0_req_0 : boolean;
  signal ptr_deref_1113_store_0_ack_0 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal ptr_deref_1113_store_0_req_1 : boolean;
  signal type_cast_1274_inst_ack_0 : boolean;
  signal ptr_deref_1113_store_0_ack_1 : boolean;
  signal type_cast_1274_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1 : boolean;
  signal W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1628_inst_ack_1 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1 : boolean;
  signal type_cast_600_inst_req_0 : boolean;
  signal W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0 : boolean;
  signal type_cast_600_inst_ack_0 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1 : boolean;
  signal W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1 : boolean;
  signal type_cast_1607_inst_req_1 : boolean;
  signal phi_stmt_1526_req_0 : boolean;
  signal type_cast_1156_inst_req_0 : boolean;
  signal type_cast_1156_inst_ack_0 : boolean;
  signal type_cast_1156_inst_req_1 : boolean;
  signal type_cast_1156_inst_ack_1 : boolean;
  signal type_cast_600_inst_req_1 : boolean;
  signal type_cast_1607_inst_ack_1 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal type_cast_1186_inst_req_1 : boolean;
  signal type_cast_1186_inst_ack_1 : boolean;
  signal type_cast_1202_inst_req_0 : boolean;
  signal type_cast_1202_inst_ack_0 : boolean;
  signal type_cast_1202_inst_req_1 : boolean;
  signal type_cast_1202_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_1 : boolean;
  signal if_stmt_1359_branch_ack_1 : boolean;
  signal if_stmt_1359_branch_ack_0 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal type_cast_1597_inst_ack_1 : boolean;
  signal call_stmt_1372_call_req_0 : boolean;
  signal call_stmt_1372_call_ack_0 : boolean;
  signal call_stmt_1372_call_req_1 : boolean;
  signal call_stmt_1372_call_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_req_1 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal type_cast_1597_inst_req_1 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_req_1 : boolean;
  signal type_cast_1385_inst_req_0 : boolean;
  signal phi_stmt_377_ack_0 : boolean;
  signal type_cast_1385_inst_ack_0 : boolean;
  signal type_cast_1385_inst_req_1 : boolean;
  signal type_cast_1385_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_ack_0 : boolean;
  signal phi_stmt_1526_ack_0 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal phi_stmt_377_req_1 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal type_cast_1395_inst_req_1 : boolean;
  signal type_cast_383_inst_ack_1 : boolean;
  signal type_cast_1395_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1622_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1637_inst_req_0 : boolean;
  signal type_cast_1405_inst_req_0 : boolean;
  signal type_cast_383_inst_req_1 : boolean;
  signal type_cast_1405_inst_ack_0 : boolean;
  signal phi_stmt_1526_req_1 : boolean;
  signal type_cast_1405_inst_req_1 : boolean;
  signal type_cast_1405_inst_ack_1 : boolean;
  signal type_cast_1532_inst_ack_1 : boolean;
  signal type_cast_1415_inst_req_0 : boolean;
  signal type_cast_383_inst_ack_0 : boolean;
  signal type_cast_1415_inst_ack_0 : boolean;
  signal type_cast_1597_inst_ack_0 : boolean;
  signal type_cast_1532_inst_req_1 : boolean;
  signal type_cast_1415_inst_req_1 : boolean;
  signal type_cast_383_inst_req_0 : boolean;
  signal type_cast_1415_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_req_1 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_ack_0 : boolean;
  signal type_cast_1532_inst_ack_0 : boolean;
  signal type_cast_1435_inst_req_0 : boolean;
  signal type_cast_1435_inst_ack_0 : boolean;
  signal type_cast_1597_inst_req_0 : boolean;
  signal type_cast_1532_inst_req_0 : boolean;
  signal type_cast_1435_inst_req_1 : boolean;
  signal type_cast_1435_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1634_inst_req_0 : boolean;
  signal type_cast_1445_inst_req_0 : boolean;
  signal type_cast_1445_inst_ack_0 : boolean;
  signal type_cast_1445_inst_req_1 : boolean;
  signal phi_stmt_377_req_0 : boolean;
  signal type_cast_1445_inst_ack_1 : boolean;
  signal phi_stmt_594_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_ack_0 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal type_cast_1455_inst_req_1 : boolean;
  signal type_cast_1455_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1619_inst_req_0 : boolean;
  signal phi_stmt_594_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1631_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1457_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1460_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1463_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1466_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1469_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1472_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1475_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1478_inst_ack_1 : boolean;
  signal if_stmt_1488_branch_req_0 : boolean;
  signal if_stmt_1488_branch_ack_1 : boolean;
  signal if_stmt_1488_branch_ack_0 : boolean;
  signal type_cast_1509_inst_req_0 : boolean;
  signal type_cast_1509_inst_ack_0 : boolean;
  signal type_cast_1509_inst_req_1 : boolean;
  signal type_cast_1509_inst_ack_1 : boolean;
  signal array_obj_ref_1538_index_offset_req_0 : boolean;
  signal array_obj_ref_1538_index_offset_ack_0 : boolean;
  signal array_obj_ref_1538_index_offset_req_1 : boolean;
  signal array_obj_ref_1538_index_offset_ack_1 : boolean;
  signal addr_of_1539_final_reg_req_0 : boolean;
  signal addr_of_1539_final_reg_ack_0 : boolean;
  signal addr_of_1539_final_reg_req_1 : boolean;
  signal addr_of_1539_final_reg_ack_1 : boolean;
  signal ptr_deref_1543_load_0_req_0 : boolean;
  signal ptr_deref_1543_load_0_ack_0 : boolean;
  signal ptr_deref_1543_load_0_req_1 : boolean;
  signal ptr_deref_1543_load_0_ack_1 : boolean;
  signal type_cast_1547_inst_req_0 : boolean;
  signal type_cast_1547_inst_ack_0 : boolean;
  signal type_cast_1547_inst_req_1 : boolean;
  signal type_cast_1547_inst_ack_1 : boolean;
  signal type_cast_1557_inst_req_0 : boolean;
  signal type_cast_1557_inst_ack_0 : boolean;
  signal type_cast_1557_inst_req_1 : boolean;
  signal type_cast_1557_inst_ack_1 : boolean;
  signal type_cast_1567_inst_req_0 : boolean;
  signal type_cast_1567_inst_ack_0 : boolean;
  signal type_cast_1567_inst_req_1 : boolean;
  signal type_cast_1567_inst_ack_1 : boolean;
  signal type_cast_1577_inst_req_0 : boolean;
  signal type_cast_1577_inst_ack_0 : boolean;
  signal type_cast_1577_inst_req_1 : boolean;
  signal type_cast_1577_inst_ack_1 : boolean;
  signal type_cast_1587_inst_req_0 : boolean;
  signal type_cast_1587_inst_ack_0 : boolean;
  signal type_cast_1587_inst_req_1 : boolean;
  signal type_cast_1587_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "concat_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  concat_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "concat_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  concat_CP_34: Block -- control-path 
    signal concat_CP_34_elements: BooleanArray(674 downto 0);
    -- 
  begin -- 
    concat_CP_34_elements(0) <= concat_CP_34_start;
    concat_CP_34_symbol <= concat_CP_34_elements(674);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (62) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_23/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/branch_block_stmt_23__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_update_start_
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Update/cr
      -- 
    rr_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => RPIPE_Concat_input_pipe_25_inst_req_0); -- 
    cr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_30_inst_req_1); -- 
    cr_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_43_inst_req_1); -- 
    cr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_55_inst_req_1); -- 
    cr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_68_inst_req_1); -- 
    cr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_80_inst_req_1); -- 
    cr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_93_inst_req_1); -- 
    cr_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_105_inst_req_1); -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_118_inst_req_1); -- 
    cr_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_130_inst_req_1); -- 
    cr_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_143_inst_req_1); -- 
    cr_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_155_inst_req_1); -- 
    cr_451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_168_inst_req_1); -- 
    cr_479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_180_inst_req_1); -- 
    cr_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_193_inst_req_1); -- 
    cr_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_205_inst_req_1); -- 
    cr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_230_inst_req_1); -- 
    cr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(0), ack => type_cast_243_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	554 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	555 
    -- CP-element group 1: 	556 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_23/do_while_stmt_817__exit__
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359__entry__
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_23/R_ifx_xend300_whilex_xend_taken_1360_place
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_1359_else_link/$entry
      -- 
    branch_req_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(1), ack => if_stmt_1359_branch_req_0); -- 
    concat_CP_34_elements(1) <= concat_CP_34_elements(554);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_update_start_
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Update/cr
      -- 
    ra_125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_0, ack => concat_CP_34_elements(2)); -- 
    cr_129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(2), ack => RPIPE_Concat_input_pipe_25_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_25_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Sample/rr
      -- 
    ca_130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_25_inst_ack_1, ack => concat_CP_34_elements(3)); -- 
    rr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(3), ack => type_cast_30_inst_req_0); -- 
    rr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(3), ack => RPIPE_Concat_input_pipe_39_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Sample/ra
      -- 
    ra_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_0, ack => concat_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	74 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_30_Update/ca
      -- 
    ca_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_30_inst_ack_1, ack => concat_CP_34_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_update_start_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Update/cr
      -- 
    ra_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_0, ack => concat_CP_34_elements(6)); -- 
    cr_157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(6), ack => RPIPE_Concat_input_pipe_39_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	10 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_39_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Sample/rr
      -- 
    ca_158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_39_inst_ack_1, ack => concat_CP_34_elements(7)); -- 
    rr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(7), ack => type_cast_43_inst_req_0); -- 
    rr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(7), ack => RPIPE_Concat_input_pipe_51_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Sample/ra
      -- 
    ra_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_0, ack => concat_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	74 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_43_Update/ca
      -- 
    ca_172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_1, ack => concat_CP_34_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_update_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Update/cr
      -- 
    ra_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_0, ack => concat_CP_34_elements(10)); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(10), ack => RPIPE_Concat_input_pipe_51_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_51_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_51_inst_ack_1, ack => concat_CP_34_elements(11)); -- 
    rr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(11), ack => type_cast_55_inst_req_0); -- 
    rr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(11), ack => RPIPE_Concat_input_pipe_64_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Sample/ra
      -- 
    ra_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_0, ack => concat_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_55_Update/ca
      -- 
    ca_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_55_inst_ack_1, ack => concat_CP_34_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_update_start_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Update/cr
      -- 
    ra_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_0, ack => concat_CP_34_elements(14)); -- 
    cr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(14), ack => RPIPE_Concat_input_pipe_64_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_64_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Sample/rr
      -- 
    ca_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_64_inst_ack_1, ack => concat_CP_34_elements(15)); -- 
    rr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(15), ack => RPIPE_Concat_input_pipe_76_inst_req_0); -- 
    rr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(15), ack => type_cast_68_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Sample/ra
      -- 
    ra_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_0, ack => concat_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	74 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_68_Update/ca
      -- 
    ca_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_1, ack => concat_CP_34_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_update_start_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Update/cr
      -- 
    ra_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_0, ack => concat_CP_34_elements(18)); -- 
    cr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(18), ack => RPIPE_Concat_input_pipe_76_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_76_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Sample/rr
      -- 
    ca_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_76_inst_ack_1, ack => concat_CP_34_elements(19)); -- 
    rr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(19), ack => RPIPE_Concat_input_pipe_89_inst_req_0); -- 
    rr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(19), ack => type_cast_80_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Sample/ra
      -- 
    ra_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_0, ack => concat_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	74 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_80_Update/ca
      -- 
    ca_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_80_inst_ack_1, ack => concat_CP_34_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_update_start_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Update/cr
      -- 
    ra_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_0, ack => concat_CP_34_elements(22)); -- 
    cr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(22), ack => RPIPE_Concat_input_pipe_89_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_89_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Sample/rr
      -- 
    ca_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_89_inst_ack_1, ack => concat_CP_34_elements(23)); -- 
    rr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(23), ack => type_cast_93_inst_req_0); -- 
    rr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(23), ack => RPIPE_Concat_input_pipe_101_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Sample/ra
      -- 
    ra_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_0, ack => concat_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	74 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_93_Update/ca
      -- 
    ca_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_1, ack => concat_CP_34_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_update_start_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Update/cr
      -- 
    ra_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_0, ack => concat_CP_34_elements(26)); -- 
    cr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(26), ack => RPIPE_Concat_input_pipe_101_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_101_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Sample/rr
      -- 
    ca_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_101_inst_ack_1, ack => concat_CP_34_elements(27)); -- 
    rr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(27), ack => RPIPE_Concat_input_pipe_114_inst_req_0); -- 
    rr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(27), ack => type_cast_105_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Sample/ra
      -- 
    ra_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_0, ack => concat_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	74 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_105_Update/ca
      -- 
    ca_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_105_inst_ack_1, ack => concat_CP_34_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_update_start_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Update/cr
      -- 
    ra_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_0, ack => concat_CP_34_elements(30)); -- 
    cr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(30), ack => RPIPE_Concat_input_pipe_114_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_114_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Sample/rr
      -- 
    ca_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_114_inst_ack_1, ack => concat_CP_34_elements(31)); -- 
    rr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(31), ack => RPIPE_Concat_input_pipe_126_inst_req_0); -- 
    rr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(31), ack => type_cast_118_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Sample/ra
      -- 
    ra_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_0, ack => concat_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	74 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_118_Update/ca
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_1, ack => concat_CP_34_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_update_start_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Update/cr
      -- 
    ra_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_0, ack => concat_CP_34_elements(34)); -- 
    cr_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(34), ack => RPIPE_Concat_input_pipe_126_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_126_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Sample/rr
      -- 
    ca_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_126_inst_ack_1, ack => concat_CP_34_elements(35)); -- 
    rr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(35), ack => RPIPE_Concat_input_pipe_139_inst_req_0); -- 
    rr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(35), ack => type_cast_130_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Sample/ra
      -- 
    ra_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_0, ack => concat_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	74 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_130_Update/ca
      -- 
    ca_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_130_inst_ack_1, ack => concat_CP_34_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_update_start_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Sample/$exit
      -- 
    ra_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_0, ack => concat_CP_34_elements(38)); -- 
    cr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(38), ack => RPIPE_Concat_input_pipe_139_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_139_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Sample/rr
      -- 
    ca_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_139_inst_ack_1, ack => concat_CP_34_elements(39)); -- 
    rr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(39), ack => type_cast_143_inst_req_0); -- 
    rr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(39), ack => RPIPE_Concat_input_pipe_151_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Sample/ra
      -- 
    ra_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_0, ack => concat_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	74 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_143_Update/ca
      -- 
    ca_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_143_inst_ack_1, ack => concat_CP_34_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_update_start_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Update/cr
      -- 
    ra_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_0, ack => concat_CP_34_elements(42)); -- 
    cr_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(42), ack => RPIPE_Concat_input_pipe_151_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_151_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Sample/rr
      -- 
    ca_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_151_inst_ack_1, ack => concat_CP_34_elements(43)); -- 
    rr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(43), ack => type_cast_155_inst_req_0); -- 
    rr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(43), ack => RPIPE_Concat_input_pipe_164_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Sample/ra
      -- 
    ra_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => concat_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	74 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_155_Update/ca
      -- 
    ca_424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => concat_CP_34_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_update_start_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Update/cr
      -- 
    ra_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_0, ack => concat_CP_34_elements(46)); -- 
    cr_437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(46), ack => RPIPE_Concat_input_pipe_164_inst_req_1); -- 
    -- CP-element group 47:  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	50 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_164_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Sample/rr
      -- 
    ca_438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_164_inst_ack_1, ack => concat_CP_34_elements(47)); -- 
    rr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(47), ack => type_cast_168_inst_req_0); -- 
    rr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(47), ack => RPIPE_Concat_input_pipe_176_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Sample/ra
      -- 
    ra_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_0, ack => concat_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	74 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_168_Update/ca
      -- 
    ca_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_168_inst_ack_1, ack => concat_CP_34_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	47 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_update_start_
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Update/cr
      -- 
    ra_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_0, ack => concat_CP_34_elements(50)); -- 
    cr_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(50), ack => RPIPE_Concat_input_pipe_176_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_176_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Sample/rr
      -- 
    ca_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_176_inst_ack_1, ack => concat_CP_34_elements(51)); -- 
    rr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(51), ack => type_cast_180_inst_req_0); -- 
    rr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(51), ack => RPIPE_Concat_input_pipe_189_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Sample/ra
      -- 
    ra_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_0, ack => concat_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	74 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_180_Update/ca
      -- 
    ca_480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_180_inst_ack_1, ack => concat_CP_34_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_update_start_
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Update/cr
      -- 
    ra_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_189_inst_ack_0, ack => concat_CP_34_elements(54)); -- 
    cr_493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(54), ack => RPIPE_Concat_input_pipe_189_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_189_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Sample/rr
      -- 
    ca_494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_189_inst_ack_1, ack => concat_CP_34_elements(55)); -- 
    rr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(55), ack => type_cast_193_inst_req_0); -- 
    rr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(55), ack => RPIPE_Concat_input_pipe_201_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Sample/ra
      -- 
    ra_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_0, ack => concat_CP_34_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	74 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_193_Update/ca
      -- 
    ca_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_193_inst_ack_1, ack => concat_CP_34_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Update/cr
      -- 
    ra_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_201_inst_ack_0, ack => concat_CP_34_elements(58)); -- 
    cr_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(58), ack => RPIPE_Concat_input_pipe_201_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_201_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Sample/rr
      -- 
    ca_522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_201_inst_ack_1, ack => concat_CP_34_elements(59)); -- 
    rr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(59), ack => type_cast_205_inst_req_0); -- 
    rr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(59), ack => RPIPE_Concat_input_pipe_214_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Sample/ra
      -- 
    ra_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => concat_CP_34_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	74 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_205_Update/ca
      -- 
    ca_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => concat_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_update_start_
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Update/cr
      -- 
    ra_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_214_inst_ack_0, ack => concat_CP_34_elements(62)); -- 
    cr_549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(62), ack => RPIPE_Concat_input_pipe_214_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_214_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Sample/rr
      -- 
    ca_550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_214_inst_ack_1, ack => concat_CP_34_elements(63)); -- 
    rr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(63), ack => type_cast_218_inst_req_0); -- 
    rr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(63), ack => RPIPE_Concat_input_pipe_226_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Sample/ra
      -- 
    ra_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => concat_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	74 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_218_Update/ca
      -- 
    ca_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => concat_CP_34_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_update_start_
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Update/cr
      -- 
    ra_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_226_inst_ack_0, ack => concat_CP_34_elements(66)); -- 
    cr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(66), ack => RPIPE_Concat_input_pipe_226_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_226_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Sample/rr
      -- 
    ca_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_226_inst_ack_1, ack => concat_CP_34_elements(67)); -- 
    rr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(67), ack => type_cast_230_inst_req_0); -- 
    rr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(67), ack => RPIPE_Concat_input_pipe_239_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Sample/ra
      -- 
    ra_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_0, ack => concat_CP_34_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_230_Update/ca
      -- 
    ca_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_230_inst_ack_1, ack => concat_CP_34_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_update_start_
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Update/cr
      -- 
    ra_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_239_inst_ack_0, ack => concat_CP_34_elements(70)); -- 
    cr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(70), ack => RPIPE_Concat_input_pipe_239_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/RPIPE_Concat_input_pipe_239_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Sample/rr
      -- 
    ca_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_239_inst_ack_1, ack => concat_CP_34_elements(71)); -- 
    rr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(71), ack => type_cast_243_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Sample/ra
      -- 
    ra_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_0, ack => concat_CP_34_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/type_cast_243_Update/ca
      -- 
    ca_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_1, ack => concat_CP_34_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	41 
    -- CP-element group 74: 	45 
    -- CP-element group 74: 	49 
    -- CP-element group 74: 	53 
    -- CP-element group 74: 	25 
    -- CP-element group 74: 	17 
    -- CP-element group 74: 	21 
    -- CP-element group 74: 	37 
    -- CP-element group 74: 	13 
    -- CP-element group 74: 	29 
    -- CP-element group 74: 	33 
    -- CP-element group 74: 	57 
    -- CP-element group 74: 	61 
    -- CP-element group 74: 	65 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	5 
    -- CP-element group 74: 	9 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307__exit__
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308__entry__
      -- CP-element group 74: 	 branch_block_stmt_23/assign_stmt_26_to_assign_stmt_307/$exit
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_23/R_cmp467_309_place
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_23/if_stmt_308_else_link/$entry
      -- 
    branch_req_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(74), ack => if_stmt_308_branch_req_0); -- 
    concat_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 17) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1);
      constant place_markings: IntegerArray(0 to 17)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant place_delays: IntegerArray(0 to 17) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 18); -- 
    begin -- 
      preds <= concat_CP_34_elements(41) & concat_CP_34_elements(45) & concat_CP_34_elements(49) & concat_CP_34_elements(53) & concat_CP_34_elements(25) & concat_CP_34_elements(17) & concat_CP_34_elements(21) & concat_CP_34_elements(37) & concat_CP_34_elements(13) & concat_CP_34_elements(29) & concat_CP_34_elements(33) & concat_CP_34_elements(57) & concat_CP_34_elements(61) & concat_CP_34_elements(65) & concat_CP_34_elements(69) & concat_CP_34_elements(73) & concat_CP_34_elements(5) & concat_CP_34_elements(9);
      gj_concat_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 18, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75:  members (18) 
      -- CP-element group 75: 	 branch_block_stmt_23/merge_stmt_329__exit__
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374__entry__
      -- CP-element group 75: 	 branch_block_stmt_23/merge_stmt_329_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_23/if_stmt_308_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_23/if_stmt_308_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_23/entry_bbx_xnph469
      -- CP-element group 75: 	 branch_block_stmt_23/entry_bbx_xnph469_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/$entry
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_update_start_
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_23/merge_stmt_329_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_23/merge_stmt_329_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_23/merge_stmt_329_PhiAck/dummy
      -- 
    if_choice_transition_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_308_branch_ack_1, ack => concat_CP_34_elements(75)); -- 
    rr_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(75), ack => type_cast_360_inst_req_0); -- 
    cr_677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(75), ack => type_cast_360_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	654 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_308_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_23/if_stmt_308_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader
      -- CP-element group 76: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_23/entry_forx_xcond171x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_308_branch_ack_0, ack => concat_CP_34_elements(76)); -- 
    -- CP-element group 77:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	654 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77:  members (18) 
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_546__exit__
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591__entry__
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_update_start_
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_23/if_stmt_323_if_link/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/if_stmt_323_if_link/if_choice_transition
      -- CP-element group 77: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465
      -- CP-element group 77: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_546_PhiReqMerge
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_546_PhiAck/dummy
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_546_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/merge_stmt_546_PhiAck/$entry
      -- CP-element group 77: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$exit
      -- CP-element group 77: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$entry
      -- 
    if_choice_transition_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_323_branch_ack_1, ack => concat_CP_34_elements(77)); -- 
    cr_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(77), ack => type_cast_577_inst_req_1); -- 
    rr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(77), ack => type_cast_577_inst_req_0); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	654 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	667 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_23/if_stmt_323_else_link/$exit
      -- CP-element group 78: 	 branch_block_stmt_23/if_stmt_323_else_link/else_choice_transition
      -- CP-element group 78: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231
      -- CP-element group 78: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_23/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$entry
      -- 
    else_choice_transition_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_323_branch_ack_0, ack => concat_CP_34_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Sample/ra
      -- 
    ra_673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_0, ack => concat_CP_34_elements(79)); -- 
    -- CP-element group 80:  transition  place  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	655 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374__exit__
      -- CP-element group 80: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/$exit
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_23/assign_stmt_334_to_assign_stmt_374/type_cast_360_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/$entry
      -- CP-element group 80: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/$entry
      -- 
    ca_678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_1, ack => concat_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	660 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	120 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_sample_complete
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Sample/ack
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_389_index_offset_ack_0, ack => concat_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	660 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (11) 
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_root_address_calculated
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_offset_calculated
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_base_plus_offset/$entry
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_base_plus_offset/$exit
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_base_plus_offset/sum_rename_req
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_base_plus_offset/sum_rename_ack
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_request/$entry
      -- CP-element group 82: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_request/req
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_389_index_offset_ack_1, ack => concat_CP_34_elements(82)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(82), ack => addr_of_390_final_reg_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_request/$exit
      -- CP-element group 83: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_request/ack
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_390_final_reg_ack_0, ack => concat_CP_34_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	660 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	117 
    -- CP-element group 84:  members (19) 
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_word_addrgen/root_register_ack
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_word_addrgen/root_register_req
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_word_addrgen/$exit
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_complete/ack
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_word_addrgen/$entry
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_plus_offset/sum_rename_ack
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_word_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_root_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_address_resized
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_addr_resize/$entry
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_addr_resize/$exit
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_addr_resize/base_resize_req
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_addr_resize/base_resize_ack
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_plus_offset/$entry
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_plus_offset/$exit
      -- CP-element group 84: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_base_plus_offset/sum_rename_req
      -- 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_390_final_reg_ack_1, ack => concat_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	660 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_update_start_
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Update/cr
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_393_inst_ack_0, ack => concat_CP_34_elements(85)); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(85), ack => RPIPE_Concat_input_pipe_393_inst_req_1); -- 
    -- CP-element group 86:  fork  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	89 
    -- CP-element group 86:  members (9) 
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Sample/rr
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_393_inst_ack_1, ack => concat_CP_34_elements(86)); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(86), ack => type_cast_397_inst_req_0); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(86), ack => RPIPE_Concat_input_pipe_406_inst_req_0); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Sample/ra
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_0, ack => concat_CP_34_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	660 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	117 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Update/ca
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_1, ack => concat_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	86 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_update_start_
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Update/cr
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_406_inst_ack_0, ack => concat_CP_34_elements(89)); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(89), ack => RPIPE_Concat_input_pipe_406_inst_req_1); -- 
    -- CP-element group 90:  fork  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	93 
    -- CP-element group 90:  members (9) 
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_406_Update/$exit
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_406_inst_ack_1, ack => concat_CP_34_elements(90)); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(90), ack => type_cast_410_inst_req_0); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(90), ack => RPIPE_Concat_input_pipe_424_inst_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_0, ack => concat_CP_34_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	660 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	117 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_1, ack => concat_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_update_start_
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Update/cr
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_424_inst_ack_0, ack => concat_CP_34_elements(93)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(93), ack => RPIPE_Concat_input_pipe_424_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	97 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_424_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Sample/rr
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_424_inst_ack_1, ack => concat_CP_34_elements(94)); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(94), ack => type_cast_428_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(94), ack => RPIPE_Concat_input_pipe_442_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_428_inst_ack_0, ack => concat_CP_34_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	660 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	117 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_428_inst_ack_1, ack => concat_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	94 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_update_start_
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_442_inst_ack_0, ack => concat_CP_34_elements(97)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(97), ack => RPIPE_Concat_input_pipe_442_inst_req_1); -- 
    -- CP-element group 98:  fork  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: 	101 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_442_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_442_inst_ack_1, ack => concat_CP_34_elements(98)); -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(98), ack => type_cast_446_inst_req_0); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(98), ack => RPIPE_Concat_input_pipe_460_inst_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Sample/ra
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_0, ack => concat_CP_34_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	660 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	117 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_446_inst_ack_1, ack => concat_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	98 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_update_start_
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Update/cr
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_460_inst_ack_0, ack => concat_CP_34_elements(101)); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(101), ack => RPIPE_Concat_input_pipe_460_inst_req_1); -- 
    -- CP-element group 102:  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	105 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_460_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Sample/rr
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_460_inst_ack_1, ack => concat_CP_34_elements(102)); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(102), ack => type_cast_464_inst_req_0); -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(102), ack => RPIPE_Concat_input_pipe_478_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Sample/ra
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_464_inst_ack_0, ack => concat_CP_34_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	660 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	117 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Update/ca
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_464_inst_ack_1, ack => concat_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_update_start_
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Update/cr
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_478_inst_ack_0, ack => concat_CP_34_elements(105)); -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(105), ack => RPIPE_Concat_input_pipe_478_inst_req_1); -- 
    -- CP-element group 106:  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_478_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Sample/rr
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_478_inst_ack_1, ack => concat_CP_34_elements(106)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(106), ack => type_cast_482_inst_req_0); -- 
    rr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(106), ack => RPIPE_Concat_input_pipe_496_inst_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_0, ack => concat_CP_34_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	660 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	117 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_482_inst_ack_1, ack => concat_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_update_start_
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Update/cr
      -- 
    ra_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_496_inst_ack_0, ack => concat_CP_34_elements(109)); -- 
    cr_908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(109), ack => RPIPE_Concat_input_pipe_496_inst_req_1); -- 
    -- CP-element group 110:  fork  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_496_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Sample/rr
      -- 
    ca_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_496_inst_ack_1, ack => concat_CP_34_elements(110)); -- 
    rr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(110), ack => type_cast_500_inst_req_0); -- 
    rr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(110), ack => RPIPE_Concat_input_pipe_514_inst_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Sample/ra
      -- 
    ra_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_0, ack => concat_CP_34_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	660 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	117 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Update/ca
      -- 
    ca_923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_500_inst_ack_1, ack => concat_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_update_start_
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Update/cr
      -- 
    ra_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_514_inst_ack_0, ack => concat_CP_34_elements(113)); -- 
    cr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(113), ack => RPIPE_Concat_input_pipe_514_inst_req_1); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_514_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Sample/rr
      -- 
    ca_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_514_inst_ack_1, ack => concat_CP_34_elements(114)); -- 
    rr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(114), ack => type_cast_518_inst_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Sample/ra
      -- 
    ra_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_0, ack => concat_CP_34_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	660 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Update/ca
      -- 
    ca_951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_518_inst_ack_1, ack => concat_CP_34_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	84 
    -- CP-element group 117: 	88 
    -- CP-element group 117: 	92 
    -- CP-element group 117: 	96 
    -- CP-element group 117: 	100 
    -- CP-element group 117: 	104 
    -- CP-element group 117: 	108 
    -- CP-element group 117: 	112 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (9) 
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/word_0/rr
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/$entry
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/ptr_deref_526_Split/split_ack
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/ptr_deref_526_Split/split_req
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/ptr_deref_526_Split/$exit
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/ptr_deref_526_Split/$entry
      -- CP-element group 117: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_sample_start_
      -- 
    rr_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(117), ack => ptr_deref_526_store_0_req_0); -- 
    concat_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(84) & concat_CP_34_elements(88) & concat_CP_34_elements(92) & concat_CP_34_elements(96) & concat_CP_34_elements(100) & concat_CP_34_elements(104) & concat_CP_34_elements(108) & concat_CP_34_elements(112) & concat_CP_34_elements(116);
      gj_concat_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/word_0/ra
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Sample/word_access_start/$exit
      -- CP-element group 118: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_sample_completed_
      -- 
    ra_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_526_store_0_ack_0, ack => concat_CP_34_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	660 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/word_0/ca
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/$exit
      -- CP-element group 119: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_update_completed_
      -- 
    ca_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_526_store_0_ack_1, ack => concat_CP_34_elements(119)); -- 
    -- CP-element group 120:  branch  join  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	81 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (10) 
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_dead_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539__exit__
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540__entry__
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_else_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/$exit
      -- CP-element group 120: 	 branch_block_stmt_23/R_exitcond2_541_place
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_if_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_23/if_stmt_540_eval_test/$entry
      -- 
    branch_req_1009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(120), ack => if_stmt_540_branch_req_0); -- 
    concat_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(81) & concat_CP_34_elements(119);
      gj_concat_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  transition  place  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	654 
    -- CP-element group 121:  members (13) 
      -- CP-element group 121: 	 branch_block_stmt_23/merge_stmt_314__exit__
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit
      -- CP-element group 121: 	 branch_block_stmt_23/if_stmt_540_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_23/if_stmt_540_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_23/merge_stmt_314_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_23/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_23/merge_stmt_314_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_23/merge_stmt_314_PhiAck/dummy
      -- CP-element group 121: 	 branch_block_stmt_23/merge_stmt_314_PhiAck/$exit
      -- 
    if_choice_transition_1014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_540_branch_ack_1, ack => concat_CP_34_elements(121)); -- 
    -- CP-element group 122:  fork  transition  place  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	656 
    -- CP-element group 122: 	657 
    -- CP-element group 122:  members (12) 
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/if_stmt_540_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody
      -- CP-element group 122: 	 branch_block_stmt_23/if_stmt_540_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Update/cr
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_540_branch_ack_0, ack => concat_CP_34_elements(122)); -- 
    cr_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(122), ack => type_cast_383_inst_req_1); -- 
    rr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(122), ack => type_cast_383_inst_req_0); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Sample/ra
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_sample_completed_
      -- 
    ra_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => concat_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	661 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591__exit__
      -- CP-element group 124: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/type_cast_577_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_23/assign_stmt_551_to_assign_stmt_591/$exit
      -- CP-element group 124: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/$entry
      -- CP-element group 124: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/$entry
      -- 
    ca_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => concat_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	666 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Sample/ack
      -- CP-element group 125: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Sample/$exit
      -- 
    ack_1066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_offset_ack_0, ack => concat_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	666 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_request/req
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Update/$exit
      -- 
    ack_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_606_index_offset_ack_1, ack => concat_CP_34_elements(126)); -- 
    req_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(126), ack => addr_of_607_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_request/ack
      -- CP-element group 127: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_request/$exit
      -- 
    ack_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_607_final_reg_ack_0, ack => concat_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	666 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_complete/ack
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_base_address_resized
      -- 
    ack_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_607_final_reg_ack_1, ack => concat_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	666 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_update_start_
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Update/cr
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_610_inst_ack_0, ack => concat_CP_34_elements(129)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(129), ack => RPIPE_Concat_input_pipe_610_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Update/$exit
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_610_inst_ack_1, ack => concat_CP_34_elements(130)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(130), ack => type_cast_614_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(130), ack => RPIPE_Concat_input_pipe_623_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Sample/$exit
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => concat_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	666 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_update_completed_
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_1, ack => concat_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_update_start_
      -- CP-element group 133: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_623_inst_ack_0, ack => concat_CP_34_elements(133)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(133), ack => RPIPE_Concat_input_pipe_623_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_623_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_sample_start_
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_623_inst_ack_1, ack => concat_CP_34_elements(134)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(134), ack => type_cast_627_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(134), ack => RPIPE_Concat_input_pipe_641_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_sample_completed_
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_0, ack => concat_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	666 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_update_completed_
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_627_inst_ack_1, ack => concat_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_update_start_
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Sample/$exit
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_641_inst_ack_0, ack => concat_CP_34_elements(137)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(137), ack => RPIPE_Concat_input_pipe_641_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_641_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_sample_start_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_641_inst_ack_1, ack => concat_CP_34_elements(138)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(138), ack => type_cast_645_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(138), ack => RPIPE_Concat_input_pipe_659_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_sample_completed_
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_0, ack => concat_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	666 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Update/$exit
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_1, ack => concat_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_update_start_
      -- CP-element group 141: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_sample_completed_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_659_inst_ack_0, ack => concat_CP_34_elements(141)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(141), ack => RPIPE_Concat_input_pipe_659_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_659_update_completed_
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_659_inst_ack_1, ack => concat_CP_34_elements(142)); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(142), ack => type_cast_663_inst_req_0); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(142), ack => RPIPE_Concat_input_pipe_677_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_sample_completed_
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_0, ack => concat_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	666 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_update_completed_
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_663_inst_ack_1, ack => concat_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_update_start_
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Sample/ra
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_677_inst_ack_0, ack => concat_CP_34_elements(145)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(145), ack => RPIPE_Concat_input_pipe_677_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_677_Update/ca
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_677_inst_ack_1, ack => concat_CP_34_elements(146)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(146), ack => type_cast_681_inst_req_0); -- 
    rr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(146), ack => RPIPE_Concat_input_pipe_695_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_sample_completed_
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_681_inst_ack_0, ack => concat_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	666 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_update_completed_
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_681_inst_ack_1, ack => concat_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_update_start_
      -- CP-element group 149: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_sample_completed_
      -- 
    ra_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_695_inst_ack_0, ack => concat_CP_34_elements(149)); -- 
    cr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(149), ack => RPIPE_Concat_input_pipe_695_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_695_Update/ca
      -- 
    ca_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_695_inst_ack_1, ack => concat_CP_34_elements(150)); -- 
    rr_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(150), ack => type_cast_699_inst_req_0); -- 
    rr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(150), ack => RPIPE_Concat_input_pipe_713_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_sample_completed_
      -- 
    ra_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => concat_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	666 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_update_completed_
      -- 
    ca_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => concat_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_update_start_
      -- 
    ra_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_713_inst_ack_0, ack => concat_CP_34_elements(153)); -- 
    cr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(153), ack => RPIPE_Concat_input_pipe_713_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_713_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Sample/$entry
      -- 
    ca_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_713_inst_ack_1, ack => concat_CP_34_elements(154)); -- 
    rr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(154), ack => type_cast_717_inst_req_0); -- 
    rr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(154), ack => RPIPE_Concat_input_pipe_731_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Sample/$exit
      -- 
    ra_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_0, ack => concat_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	666 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Update/$exit
      -- 
    ca_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_1, ack => concat_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_update_start_
      -- CP-element group 157: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_sample_completed_
      -- 
    ra_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_731_inst_ack_0, ack => concat_CP_34_elements(157)); -- 
    cr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(157), ack => RPIPE_Concat_input_pipe_731_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_731_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_sample_start_
      -- 
    ca_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_731_inst_ack_1, ack => concat_CP_34_elements(158)); -- 
    rr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(158), ack => type_cast_735_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_sample_completed_
      -- 
    ra_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_0, ack => concat_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	666 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_update_completed_
      -- 
    ca_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_1, ack => concat_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/ptr_deref_743_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/ptr_deref_743_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/ptr_deref_743_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/ptr_deref_743_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/$entry
      -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(161), ack => ptr_deref_743_store_0_req_0); -- 
    concat_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(128) & concat_CP_34_elements(132) & concat_CP_34_elements(136) & concat_CP_34_elements(140) & concat_CP_34_elements(144) & concat_CP_34_elements(148) & concat_CP_34_elements(152) & concat_CP_34_elements(156) & concat_CP_34_elements(160);
      gj_concat_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Sample/$exit
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_store_0_ack_0, ack => concat_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	666 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/word_0/ca
      -- 
    ca_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_store_0_ack_1, ack => concat_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	125 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756__exit__
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757__entry__
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/$exit
      -- CP-element group 164: 	 branch_block_stmt_23/R_exitcond_758_place
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_23/if_stmt_757_dead_link/$entry
      -- 
    branch_req_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(164), ack => if_stmt_757_branch_req_0); -- 
    concat_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(125) & concat_CP_34_elements(163);
      gj_concat_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	667 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_23/merge_stmt_763__exit__
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231
      -- CP-element group 165: 	 branch_block_stmt_23/if_stmt_757_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_23/if_stmt_757_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_23/merge_stmt_763_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xend231x_xloopexit_forx_xend231_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/merge_stmt_763_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_23/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_757_branch_ack_1, ack => concat_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	662 
    -- CP-element group 166: 	663 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/if_stmt_757_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_23/if_stmt_757_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_757_branch_ack_0, ack => concat_CP_34_elements(166)); -- 
    rr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(166), ack => type_cast_600_inst_req_0); -- 
    cr_3600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(166), ack => type_cast_600_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	667 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/cra
      -- CP-element group 167: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/$exit
      -- 
    cra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_768_call_ack_0, ack => concat_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	667 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (17) 
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787/$exit
      -- CP-element group 168: 	 branch_block_stmt_23/call_stmt_768/$exit
      -- CP-element group 168: 	 branch_block_stmt_23/call_stmt_768__exit__
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787__entry__
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787__exit__
      -- CP-element group 168: 	 branch_block_stmt_23/forx_xend231_whilex_xbody
      -- CP-element group 168: 	 branch_block_stmt_23/merge_stmt_789__exit__
      -- CP-element group 168: 	 branch_block_stmt_23/do_while_stmt_817__entry__
      -- CP-element group 168: 	 branch_block_stmt_23/assign_stmt_775_to_assign_stmt_787/$entry
      -- CP-element group 168: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/cca
      -- CP-element group 168: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_23/merge_stmt_789_PhiAck/$exit
      -- CP-element group 168: 	 branch_block_stmt_23/merge_stmt_789_PhiAck/$entry
      -- CP-element group 168: 	 branch_block_stmt_23/merge_stmt_789_PhiReqMerge
      -- CP-element group 168: 	 branch_block_stmt_23/forx_xend231_whilex_xbody_PhiReq/$exit
      -- CP-element group 168: 	 branch_block_stmt_23/forx_xend231_whilex_xbody_PhiReq/$entry
      -- 
    cca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_768_call_ack_1, ack => concat_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  place  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	175 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817__entry__
      -- CP-element group 169: 	 branch_block_stmt_23/do_while_stmt_817/$entry
      -- 
    concat_CP_34_elements(169) <= concat_CP_34_elements(168);
    -- CP-element group 170:  merge  place  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	554 
    -- CP-element group 170:  members (1) 
      -- CP-element group 170: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817__exit__
      -- 
    -- Element group concat_CP_34_elements(170) is bound as output of CP function.
    -- CP-element group 171:  merge  place  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	174 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_23/do_while_stmt_817/loop_back
      -- 
    -- Element group concat_CP_34_elements(171) is bound as output of CP function.
    -- CP-element group 172:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	177 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	552 
    -- CP-element group 172: 	553 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_817/condition_done
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/$entry
      -- CP-element group 172: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/$entry
      -- 
    concat_CP_34_elements(172) <= concat_CP_34_elements(177);
    -- CP-element group 173:  branch  place  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	551 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_23/do_while_stmt_817/loop_body_done
      -- 
    concat_CP_34_elements(173) <= concat_CP_34_elements(551);
    -- CP-element group 174:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	171 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	186 
    -- CP-element group 174: 	207 
    -- CP-element group 174: 	228 
    -- CP-element group 174: 	249 
    -- CP-element group 174: 	270 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/back_edge_to_loop_body
      -- 
    concat_CP_34_elements(174) <= concat_CP_34_elements(171);
    -- CP-element group 175:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	169 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	188 
    -- CP-element group 175: 	209 
    -- CP-element group 175: 	230 
    -- CP-element group 175: 	251 
    -- CP-element group 175: 	272 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/first_time_through_loop_body
      -- 
    concat_CP_34_elements(175) <= concat_CP_34_elements(169);
    -- CP-element group 176:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	182 
    -- CP-element group 176: 	183 
    -- CP-element group 176: 	201 
    -- CP-element group 176: 	202 
    -- CP-element group 176: 	222 
    -- CP-element group 176: 	223 
    -- CP-element group 176: 	243 
    -- CP-element group 176: 	244 
    -- CP-element group 176: 	264 
    -- CP-element group 176: 	265 
    -- CP-element group 176: 	298 
    -- CP-element group 176: 	299 
    -- CP-element group 176: 	321 
    -- CP-element group 176: 	322 
    -- CP-element group 176: 	408 
    -- CP-element group 176: 	409 
    -- CP-element group 176: 	431 
    -- CP-element group 176: 	432 
    -- CP-element group 176: 	549 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/loop_body_start
      -- CP-element group 176: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/$entry
      -- 
    -- Element group concat_CP_34_elements(176) is bound as output of CP function.
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	181 
    -- CP-element group 177: 	548 
    -- CP-element group 177: 	549 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	172 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/condition_evaluated
      -- 
    condition_evaluated_1414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(177), ack => do_while_stmt_817_branch_req_0); -- 
    concat_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(181) & concat_CP_34_elements(548) & concat_CP_34_elements(549);
      gj_concat_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	182 
    -- CP-element group 178: 	201 
    -- CP-element group 178: 	222 
    -- CP-element group 178: 	243 
    -- CP-element group 178: 	264 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	181 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178: 	224 
    -- CP-element group 178: 	245 
    -- CP-element group 178: 	266 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_sample_req
      -- CP-element group 178: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_start__ps
      -- 
    concat_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(182) & concat_CP_34_elements(201) & concat_CP_34_elements(222) & concat_CP_34_elements(243) & concat_CP_34_elements(264) & concat_CP_34_elements(181);
      gj_concat_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	184 
    -- CP-element group 179: 	204 
    -- CP-element group 179: 	225 
    -- CP-element group 179: 	246 
    -- CP-element group 179: 	267 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	286 
    -- CP-element group 179: 	344 
    -- CP-element group 179: 	356 
    -- CP-element group 179: 	474 
    -- CP-element group 179: 	482 
    -- CP-element group 179: 	486 
    -- CP-element group 179: 	490 
    -- CP-element group 179: 	494 
    -- CP-element group 179: 	502 
    -- CP-element group 179: 	506 
    -- CP-element group 179: 	510 
    -- CP-element group 179: 	518 
    -- CP-element group 179: 	522 
    -- CP-element group 179: 	530 
    -- CP-element group 179: 	534 
    -- CP-element group 179: 	542 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	182 
    -- CP-element group 179: 	201 
    -- CP-element group 179: 	222 
    -- CP-element group 179: 	243 
    -- CP-element group 179: 	264 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_sample_ack
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_completed_
      -- 
    concat_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(184) & concat_CP_34_elements(204) & concat_CP_34_elements(225) & concat_CP_34_elements(246) & concat_CP_34_elements(267);
      gj_concat_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	183 
    -- CP-element group 180: 	202 
    -- CP-element group 180: 	223 
    -- CP-element group 180: 	244 
    -- CP-element group 180: 	265 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180: 	226 
    -- CP-element group 180: 	247 
    -- CP-element group 180: 	268 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_start__ps
      -- CP-element group 180: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_update_req
      -- 
    concat_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(183) & concat_CP_34_elements(202) & concat_CP_34_elements(223) & concat_CP_34_elements(244) & concat_CP_34_elements(265);
      gj_concat_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	185 
    -- CP-element group 181: 	206 
    -- CP-element group 181: 	227 
    -- CP-element group 181: 	248 
    -- CP-element group 181: 	269 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	177 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	178 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/aggregated_phi_update_ack
      -- 
    concat_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(185) & concat_CP_34_elements(206) & concat_CP_34_elements(227) & concat_CP_34_elements(248) & concat_CP_34_elements(269);
      gj_concat_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	176 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: 	476 
    -- CP-element group 182: 	484 
    -- CP-element group 182: 	488 
    -- CP-element group 182: 	508 
    -- CP-element group 182: 	512 
    -- CP-element group 182: 	520 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	178 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_start_
      -- 
    concat_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(179) & concat_CP_34_elements(476) & concat_CP_34_elements(484) & concat_CP_34_elements(488) & concat_CP_34_elements(508) & concat_CP_34_elements(512) & concat_CP_34_elements(520);
      gj_concat_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	176 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: 	314 
    -- CP-element group 183: 	349 
    -- CP-element group 183: 	353 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	180 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_start_
      -- 
    concat_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(185) & concat_CP_34_elements(314) & concat_CP_34_elements(349) & concat_CP_34_elements(353);
      gj_concat_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	179 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(184) is bound as output of CP function.
    -- CP-element group 185:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	181 
    -- CP-element group 185: 	312 
    -- CP-element group 185: 	347 
    -- CP-element group 185: 	351 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	183 
    -- CP-element group 185:  members (2) 
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_completed__ps
      -- CP-element group 185: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_update_completed_
      -- 
    -- Element group concat_CP_34_elements(185) is bound as output of CP function.
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	174 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_trigger
      -- 
    concat_CP_34_elements(186) <= concat_CP_34_elements(174);
    -- CP-element group 187:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (2) 
      -- CP-element group 187: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_sample_req
      -- CP-element group 187: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_loopback_sample_req_ps
      -- 
    phi_stmt_819_loopback_sample_req_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_819_loopback_sample_req_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(187), ack => phi_stmt_819_req_0); -- 
    -- Element group concat_CP_34_elements(187) is bound as output of CP function.
    -- CP-element group 188:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	175 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_trigger
      -- 
    concat_CP_34_elements(188) <= concat_CP_34_elements(175);
    -- CP-element group 189:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_sample_req
      -- CP-element group 189: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_entry_sample_req_ps
      -- 
    phi_stmt_819_entry_sample_req_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_819_entry_sample_req_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(189), ack => phi_stmt_819_req_1); -- 
    -- Element group concat_CP_34_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (2) 
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_phi_mux_ack
      -- CP-element group 190: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_819_phi_mux_ack_ps
      -- 
    phi_stmt_819_phi_mux_ack_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_819_ack_0, ack => concat_CP_34_elements(190)); -- 
    -- CP-element group 191:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(191) is bound as output of CP function.
    -- CP-element group 192:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(192) is bound as output of CP function.
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/rr
      -- 
    rr_1448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(193), ack => type_cast_822_inst_req_0); -- 
    concat_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(191) & concat_CP_34_elements(195);
      gj_concat_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_start_
      -- CP-element group 194: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/cr
      -- 
    cr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(194), ack => type_cast_822_inst_req_1); -- 
    concat_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(192) & concat_CP_34_elements(196);
      gj_concat_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Sample/ra
      -- 
    ra_1449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => concat_CP_34_elements(195)); -- 
    -- CP-element group 196:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_completed__ps
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_822_Update/ca
      -- 
    ca_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => concat_CP_34_elements(196)); -- 
    -- CP-element group 197:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (4) 
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_start__ps
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_completed__ps
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(197) is bound as output of CP function.
    -- CP-element group 198:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (2) 
      -- CP-element group 198: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_start__ps
      -- CP-element group 198: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_start_
      -- 
    -- Element group concat_CP_34_elements(198) is bound as output of CP function.
    -- CP-element group 199:  join  transition  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_completed__ps
      -- 
    concat_CP_34_elements(199) <= concat_CP_34_elements(200);
    -- CP-element group 200:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	199 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_outx_x1_at_entry_823_update_completed_
      -- 
    -- Element group concat_CP_34_elements(200) is a control-delay.
    cp_element_200_delay: control_delay_element  generic map(name => " 200_delay", delay_value => 1)  port map(req => concat_CP_34_elements(198), ack => concat_CP_34_elements(200), clk => clk, reset =>reset);
    -- CP-element group 201:  join  transition  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	176 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	179 
    -- CP-element group 201: 	288 
    -- CP-element group 201: 	346 
    -- CP-element group 201: 	358 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	178 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_start_
      -- 
    concat_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(179) & concat_CP_34_elements(288) & concat_CP_34_elements(346) & concat_CP_34_elements(358);
      gj_concat_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  join  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	176 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	206 
    -- CP-element group 202: 	291 
    -- CP-element group 202: 	345 
    -- CP-element group 202: 	357 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	180 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_start_
      -- 
    concat_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(206) & concat_CP_34_elements(291) & concat_CP_34_elements(345) & concat_CP_34_elements(357);
      gj_concat_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	178 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_start__ps
      -- 
    concat_CP_34_elements(203) <= concat_CP_34_elements(178);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	179 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(204) is bound as output of CP function.
    -- CP-element group 205:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	180 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_start__ps
      -- 
    concat_CP_34_elements(205) <= concat_CP_34_elements(180);
    -- CP-element group 206:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	181 
    -- CP-element group 206: 	289 
    -- CP-element group 206: 	343 
    -- CP-element group 206: 	355 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	202 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(206) is bound as output of CP function.
    -- CP-element group 207:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_trigger
      -- 
    concat_CP_34_elements(207) <= concat_CP_34_elements(174);
    -- CP-element group 208:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_sample_req
      -- CP-element group 208: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_loopback_sample_req_ps
      -- 
    phi_stmt_824_loopback_sample_req_1473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_824_loopback_sample_req_1473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(208), ack => phi_stmt_824_req_0); -- 
    -- Element group concat_CP_34_elements(208) is bound as output of CP function.
    -- CP-element group 209:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	175 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_trigger
      -- 
    concat_CP_34_elements(209) <= concat_CP_34_elements(175);
    -- CP-element group 210:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_sample_req
      -- CP-element group 210: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_entry_sample_req_ps
      -- 
    phi_stmt_824_entry_sample_req_1476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_824_entry_sample_req_1476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(210), ack => phi_stmt_824_req_1); -- 
    -- Element group concat_CP_34_elements(210) is bound as output of CP function.
    -- CP-element group 211:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (2) 
      -- CP-element group 211: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_phi_mux_ack
      -- CP-element group 211: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_824_phi_mux_ack_ps
      -- 
    phi_stmt_824_phi_mux_ack_1479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_824_ack_0, ack => concat_CP_34_elements(211)); -- 
    -- CP-element group 212:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(212) is bound as output of CP function.
    -- CP-element group 213:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(213) is bound as output of CP function.
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/rr
      -- 
    rr_1492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(214), ack => type_cast_827_inst_req_0); -- 
    concat_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(212) & concat_CP_34_elements(216);
      gj_concat_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	217 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_start_
      -- CP-element group 215: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/cr
      -- 
    cr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(215), ack => type_cast_827_inst_req_1); -- 
    concat_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(213) & concat_CP_34_elements(217);
      gj_concat_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (4) 
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_completed__ps
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Sample/ra
      -- 
    ra_1493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_0, ack => concat_CP_34_elements(216)); -- 
    -- CP-element group 217:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: marked-successors 
    -- CP-element group 217: 	215 
    -- CP-element group 217:  members (4) 
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_completed__ps
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_827_Update/ca
      -- 
    ca_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_1, ack => concat_CP_34_elements(217)); -- 
    -- CP-element group 218:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (4) 
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_start__ps
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_completed__ps
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(218) is bound as output of CP function.
    -- CP-element group 219:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (2) 
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_start__ps
      -- CP-element group 219: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_start_
      -- 
    -- Element group concat_CP_34_elements(219) is bound as output of CP function.
    -- CP-element group 220:  join  transition  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	221 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_completed__ps
      -- 
    concat_CP_34_elements(220) <= concat_CP_34_elements(221);
    -- CP-element group 221:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	220 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp1x_x1_at_entry_828_update_completed_
      -- 
    -- Element group concat_CP_34_elements(221) is a control-delay.
    cp_element_221_delay: control_delay_element  generic map(name => " 221_delay", delay_value => 1)  port map(req => concat_CP_34_elements(219), ack => concat_CP_34_elements(221), clk => clk, reset =>reset);
    -- CP-element group 222:  join  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	176 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	179 
    -- CP-element group 222: 	476 
    -- CP-element group 222: 	484 
    -- CP-element group 222: 	488 
    -- CP-element group 222: 	492 
    -- CP-element group 222: 	496 
    -- CP-element group 222: 	504 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	178 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_start_
      -- 
    concat_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(179) & concat_CP_34_elements(476) & concat_CP_34_elements(484) & concat_CP_34_elements(488) & concat_CP_34_elements(492) & concat_CP_34_elements(496) & concat_CP_34_elements(504);
      gj_concat_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	176 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	227 
    -- CP-element group 223: 	401 
    -- CP-element group 223: 	455 
    -- CP-element group 223: 	467 
    -- CP-element group 223: 	499 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	180 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_start_
      -- 
    concat_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(227) & concat_CP_34_elements(401) & concat_CP_34_elements(455) & concat_CP_34_elements(467) & concat_CP_34_elements(499);
      gj_concat_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	178 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_start__ps
      -- 
    concat_CP_34_elements(224) <= concat_CP_34_elements(178);
    -- CP-element group 225:  join  transition  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	179 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(225) is bound as output of CP function.
    -- CP-element group 226:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	180 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_start__ps
      -- 
    concat_CP_34_elements(226) <= concat_CP_34_elements(180);
    -- CP-element group 227:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	181 
    -- CP-element group 227: 	399 
    -- CP-element group 227: 	453 
    -- CP-element group 227: 	465 
    -- CP-element group 227: 	497 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	223 
    -- CP-element group 227:  members (2) 
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(227) is bound as output of CP function.
    -- CP-element group 228:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	174 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_trigger
      -- 
    concat_CP_34_elements(228) <= concat_CP_34_elements(174);
    -- CP-element group 229:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_sample_req
      -- CP-element group 229: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_loopback_sample_req_ps
      -- 
    phi_stmt_829_loopback_sample_req_1517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_loopback_sample_req_1517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(229), ack => phi_stmt_829_req_0); -- 
    -- Element group concat_CP_34_elements(229) is bound as output of CP function.
    -- CP-element group 230:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	175 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_trigger
      -- 
    concat_CP_34_elements(230) <= concat_CP_34_elements(175);
    -- CP-element group 231:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_sample_req
      -- CP-element group 231: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_entry_sample_req_ps
      -- 
    phi_stmt_829_entry_sample_req_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_829_entry_sample_req_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(231), ack => phi_stmt_829_req_1); -- 
    -- Element group concat_CP_34_elements(231) is bound as output of CP function.
    -- CP-element group 232:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (2) 
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_phi_mux_ack
      -- CP-element group 232: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_829_phi_mux_ack_ps
      -- 
    phi_stmt_829_phi_mux_ack_1523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_829_ack_0, ack => concat_CP_34_elements(232)); -- 
    -- CP-element group 233:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(233) is bound as output of CP function.
    -- CP-element group 234:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(234) is bound as output of CP function.
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	237 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/rr
      -- 
    rr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(235), ack => type_cast_832_inst_req_0); -- 
    concat_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(233) & concat_CP_34_elements(237);
      gj_concat_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_start_
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/$entry
      -- CP-element group 236: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/cr
      -- 
    cr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(236), ack => type_cast_832_inst_req_1); -- 
    concat_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(234) & concat_CP_34_elements(238);
      gj_concat_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: marked-successors 
    -- CP-element group 237: 	235 
    -- CP-element group 237:  members (4) 
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_completed__ps
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Sample/ra
      -- 
    ra_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => concat_CP_34_elements(237)); -- 
    -- CP-element group 238:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (4) 
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_completed__ps
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_832_Update/ca
      -- 
    ca_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => concat_CP_34_elements(238)); -- 
    -- CP-element group 239:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (4) 
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_start__ps
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_completed__ps
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_start__ps
      -- CP-element group 240: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_start_
      -- 
    -- Element group concat_CP_34_elements(240) is bound as output of CP function.
    -- CP-element group 241:  join  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	242 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_completed__ps
      -- 
    concat_CP_34_elements(241) <= concat_CP_34_elements(242);
    -- CP-element group 242:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	241 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_add_inp2x_x1_at_entry_833_update_completed_
      -- 
    -- Element group concat_CP_34_elements(242) is a control-delay.
    cp_element_242_delay: control_delay_element  generic map(name => " 242_delay", delay_value => 1)  port map(req => concat_CP_34_elements(240), ack => concat_CP_34_elements(242), clk => clk, reset =>reset);
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	176 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	179 
    -- CP-element group 243: 	476 
    -- CP-element group 243: 	484 
    -- CP-element group 243: 	488 
    -- CP-element group 243: 	524 
    -- CP-element group 243: 	532 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	178 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_start_
      -- 
    concat_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(179) & concat_CP_34_elements(476) & concat_CP_34_elements(484) & concat_CP_34_elements(488) & concat_CP_34_elements(524) & concat_CP_34_elements(532);
      gj_concat_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  join  transition  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	176 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	248 
    -- CP-element group 244: 	287 
    -- CP-element group 244: 	341 
    -- CP-element group 244: 	361 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	180 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_start_
      -- 
    concat_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(248) & concat_CP_34_elements(287) & concat_CP_34_elements(341) & concat_CP_34_elements(361);
      gj_concat_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	178 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (1) 
      -- CP-element group 245: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_start__ps
      -- 
    concat_CP_34_elements(245) <= concat_CP_34_elements(178);
    -- CP-element group 246:  join  transition  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	179 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(246) is bound as output of CP function.
    -- CP-element group 247:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	180 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_start__ps
      -- 
    concat_CP_34_elements(247) <= concat_CP_34_elements(180);
    -- CP-element group 248:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	181 
    -- CP-element group 248: 	285 
    -- CP-element group 248: 	339 
    -- CP-element group 248: 	359 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	244 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(248) is bound as output of CP function.
    -- CP-element group 249:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	174 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (1) 
      -- CP-element group 249: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_trigger
      -- 
    concat_CP_34_elements(249) <= concat_CP_34_elements(174);
    -- CP-element group 250:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_sample_req
      -- CP-element group 250: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_loopback_sample_req_ps
      -- 
    phi_stmt_834_loopback_sample_req_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_834_loopback_sample_req_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(250), ack => phi_stmt_834_req_0); -- 
    -- Element group concat_CP_34_elements(250) is bound as output of CP function.
    -- CP-element group 251:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	175 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (1) 
      -- CP-element group 251: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_trigger
      -- 
    concat_CP_34_elements(251) <= concat_CP_34_elements(175);
    -- CP-element group 252:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (2) 
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_sample_req
      -- CP-element group 252: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_entry_sample_req_ps
      -- 
    phi_stmt_834_entry_sample_req_1564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_834_entry_sample_req_1564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(252), ack => phi_stmt_834_req_1); -- 
    -- Element group concat_CP_34_elements(252) is bound as output of CP function.
    -- CP-element group 253:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (2) 
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_phi_mux_ack_ps
      -- CP-element group 253: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_834_phi_mux_ack
      -- 
    phi_stmt_834_phi_mux_ack_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_834_ack_0, ack => concat_CP_34_elements(253)); -- 
    -- CP-element group 254:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (1) 
      -- CP-element group 254: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(254) is bound as output of CP function.
    -- CP-element group 255:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(255) is bound as output of CP function.
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/rr
      -- 
    rr_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(256), ack => type_cast_837_inst_req_0); -- 
    concat_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(254) & concat_CP_34_elements(258);
      gj_concat_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_start_
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/cr
      -- 
    cr_1585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(257), ack => type_cast_837_inst_req_1); -- 
    concat_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(255) & concat_CP_34_elements(259);
      gj_concat_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (4) 
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_completed__ps
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Sample/ra
      -- 
    ra_1581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => concat_CP_34_elements(258)); -- 
    -- CP-element group 259:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (4) 
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_completed__ps
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_837_Update/ca
      -- 
    ca_1586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_1, ack => concat_CP_34_elements(259)); -- 
    -- CP-element group 260:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (4) 
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_start__ps
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_completed__ps
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(260) is bound as output of CP function.
    -- CP-element group 261:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_start__ps
      -- CP-element group 261: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_start_
      -- 
    -- Element group concat_CP_34_elements(261) is bound as output of CP function.
    -- CP-element group 262:  join  transition  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	263 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_completed__ps
      -- 
    concat_CP_34_elements(262) <= concat_CP_34_elements(263);
    -- CP-element group 263:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	262 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp1x_x1_at_entry_838_update_completed_
      -- 
    -- Element group concat_CP_34_elements(263) is a control-delay.
    cp_element_263_delay: control_delay_element  generic map(name => " 263_delay", delay_value => 1)  port map(req => concat_CP_34_elements(261), ack => concat_CP_34_elements(263), clk => clk, reset =>reset);
    -- CP-element group 264:  join  transition  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	176 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	179 
    -- CP-element group 264: 	476 
    -- CP-element group 264: 	484 
    -- CP-element group 264: 	488 
    -- CP-element group 264: 	536 
    -- CP-element group 264: 	544 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	178 
    -- CP-element group 264:  members (1) 
      -- CP-element group 264: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_start_
      -- 
    concat_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(179) & concat_CP_34_elements(476) & concat_CP_34_elements(484) & concat_CP_34_elements(488) & concat_CP_34_elements(536) & concat_CP_34_elements(544);
      gj_concat_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	176 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	269 
    -- CP-element group 265: 	381 
    -- CP-element group 265: 	451 
    -- CP-element group 265: 	471 
    -- CP-element group 265: 	539 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	180 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_start_
      -- 
    concat_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(269) & concat_CP_34_elements(381) & concat_CP_34_elements(451) & concat_CP_34_elements(471) & concat_CP_34_elements(539);
      gj_concat_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	178 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (1) 
      -- CP-element group 266: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_start__ps
      -- 
    concat_CP_34_elements(266) <= concat_CP_34_elements(178);
    -- CP-element group 267:  join  transition  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	179 
    -- CP-element group 267:  members (1) 
      -- CP-element group 267: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_sample_completed__ps
      -- 
    -- Element group concat_CP_34_elements(267) is bound as output of CP function.
    -- CP-element group 268:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	180 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (1) 
      -- CP-element group 268: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_start__ps
      -- 
    concat_CP_34_elements(268) <= concat_CP_34_elements(180);
    -- CP-element group 269:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	181 
    -- CP-element group 269: 	379 
    -- CP-element group 269: 	449 
    -- CP-element group 269: 	469 
    -- CP-element group 269: 	537 
    -- CP-element group 269: marked-successors 
    -- CP-element group 269: 	265 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_update_completed__ps
      -- 
    -- Element group concat_CP_34_elements(269) is bound as output of CP function.
    -- CP-element group 270:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	174 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (1) 
      -- CP-element group 270: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_trigger
      -- 
    concat_CP_34_elements(270) <= concat_CP_34_elements(174);
    -- CP-element group 271:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_sample_req
      -- CP-element group 271: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_loopback_sample_req_ps
      -- 
    phi_stmt_839_loopback_sample_req_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_839_loopback_sample_req_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(271), ack => phi_stmt_839_req_0); -- 
    -- Element group concat_CP_34_elements(271) is bound as output of CP function.
    -- CP-element group 272:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	175 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (1) 
      -- CP-element group 272: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_trigger
      -- 
    concat_CP_34_elements(272) <= concat_CP_34_elements(175);
    -- CP-element group 273:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_sample_req
      -- CP-element group 273: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_entry_sample_req_ps
      -- 
    phi_stmt_839_entry_sample_req_1608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_839_entry_sample_req_1608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(273), ack => phi_stmt_839_req_1); -- 
    -- Element group concat_CP_34_elements(273) is bound as output of CP function.
    -- CP-element group 274:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_phi_mux_ack
      -- CP-element group 274: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/phi_stmt_839_phi_mux_ack_ps
      -- 
    phi_stmt_839_phi_mux_ack_1611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_839_ack_0, ack => concat_CP_34_elements(274)); -- 
    -- CP-element group 275:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_start__ps
      -- 
    -- Element group concat_CP_34_elements(275) is bound as output of CP function.
    -- CP-element group 276:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (1) 
      -- CP-element group 276: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_start__ps
      -- 
    -- Element group concat_CP_34_elements(276) is bound as output of CP function.
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/rr
      -- 
    rr_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(277), ack => type_cast_842_inst_req_0); -- 
    concat_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(275) & concat_CP_34_elements(279);
      gj_concat_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_start_
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/cr
      -- 
    cr_1629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(278), ack => type_cast_842_inst_req_1); -- 
    concat_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(276) & concat_CP_34_elements(280);
      gj_concat_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (4) 
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_completed__ps
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Sample/ra
      -- 
    ra_1625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => concat_CP_34_elements(279)); -- 
    -- CP-element group 280:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (4) 
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_completed__ps
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_842_Update/ca
      -- 
    ca_1630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => concat_CP_34_elements(280)); -- 
    -- CP-element group 281:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (4) 
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_start__ps
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_completed__ps
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_sample_completed_
      -- 
    -- Element group concat_CP_34_elements(281) is bound as output of CP function.
    -- CP-element group 282:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_start__ps
      -- CP-element group 282: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_start_
      -- 
    -- Element group concat_CP_34_elements(282) is bound as output of CP function.
    -- CP-element group 283:  join  transition  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	284 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_completed__ps
      -- 
    concat_CP_34_elements(283) <= concat_CP_34_elements(284);
    -- CP-element group 284:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	283 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/R_count_inp2x_x1_at_entry_843_update_completed_
      -- 
    -- Element group concat_CP_34_elements(284) is a control-delay.
    cp_element_284_delay: control_delay_element  generic map(name => " 284_delay", delay_value => 1)  port map(req => concat_CP_34_elements(282), ack => concat_CP_34_elements(284), clk => clk, reset =>reset);
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	248 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/rr
      -- 
    rr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(285), ack => type_cast_847_inst_req_0); -- 
    concat_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(248) & concat_CP_34_elements(287);
      gj_concat_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	179 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: 	295 
    -- CP-element group 286: 	306 
    -- CP-element group 286: 	318 
    -- CP-element group 286: 	329 
    -- CP-element group 286: 	365 
    -- CP-element group 286: 	369 
    -- CP-element group 286: 	373 
    -- CP-element group 286: 	377 
    -- CP-element group 286: 	424 
    -- CP-element group 286: 	459 
    -- CP-element group 286: 	463 
    -- CP-element group 286: 	515 
    -- CP-element group 286: 	523 
    -- CP-element group 286: 	527 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_update_start_
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/cr
      -- 
    cr_1652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(286), ack => type_cast_847_inst_req_1); -- 
    concat_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(288) & concat_CP_34_elements(295) & concat_CP_34_elements(306) & concat_CP_34_elements(318) & concat_CP_34_elements(329) & concat_CP_34_elements(365) & concat_CP_34_elements(369) & concat_CP_34_elements(373) & concat_CP_34_elements(377) & concat_CP_34_elements(424) & concat_CP_34_elements(459) & concat_CP_34_elements(463) & concat_CP_34_elements(515) & concat_CP_34_elements(523) & concat_CP_34_elements(527);
      gj_concat_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	244 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Sample/ra
      -- 
    ra_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => concat_CP_34_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	293 
    -- CP-element group 288: 	304 
    -- CP-element group 288: 	316 
    -- CP-element group 288: 	327 
    -- CP-element group 288: 	363 
    -- CP-element group 288: 	367 
    -- CP-element group 288: 	371 
    -- CP-element group 288: 	375 
    -- CP-element group 288: 	422 
    -- CP-element group 288: 	457 
    -- CP-element group 288: 	461 
    -- CP-element group 288: 	513 
    -- CP-element group 288: 	521 
    -- CP-element group 288: 	525 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	201 
    -- CP-element group 288: 	286 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_847_Update/ca
      -- 
    ca_1653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => concat_CP_34_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	206 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/req
      -- 
    req_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(289), ack => W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0); -- 
    concat_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(206) & concat_CP_34_elements(291);
      gj_concat_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	295 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_update_start_
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/req
      -- 
    req_1666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(290), ack => W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1); -- 
    concat_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(292) & concat_CP_34_elements(295);
      gj_concat_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	202 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Sample/ack
      -- 
    ack_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0, ack => concat_CP_34_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_866_Update/ack
      -- 
    ack_1667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1, ack => concat_CP_34_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	288 
    -- CP-element group 293: 	292 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/rr
      -- 
    rr_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(293), ack => type_cast_870_inst_req_0); -- 
    concat_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(292) & concat_CP_34_elements(295);
      gj_concat_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: 	300 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_update_start_
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/cr
      -- 
    cr_1680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(294), ack => type_cast_870_inst_req_1); -- 
    concat_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(296) & concat_CP_34_elements(300);
      gj_concat_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	286 
    -- CP-element group 295: 	290 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Sample/ra
      -- 
    ra_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_0, ack => concat_CP_34_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	300 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (16) 
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_870_Update/ca
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resized_1
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scaled_1
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_computed_1
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/index_resize_req
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_resize_1/index_resize_ack
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/$exit
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/scale_rename_req
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_index_scale_1/scale_rename_ack
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/req
      -- 
    ca_1681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_1, ack => concat_CP_34_elements(296)); -- 
    req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(296), ack => array_obj_ref_876_index_offset_req_0); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	301 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	302 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	302 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/$entry
      -- CP-element group 297: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/req
      -- 
    req_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(297), ack => addr_of_877_final_reg_req_0); -- 
    concat_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(301) & concat_CP_34_elements(302);
      gj_concat_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	176 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	303 
    -- CP-element group 298: 	310 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	303 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_update_start_
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/$entry
      -- CP-element group 298: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/req
      -- 
    req_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(298), ack => addr_of_877_final_reg_req_1); -- 
    concat_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(303) & concat_CP_34_elements(310);
      gj_concat_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	176 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	301 
    -- CP-element group 299: 	302 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_update_start
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/req
      -- 
    req_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(299), ack => array_obj_ref_876_index_offset_req_1); -- 
    concat_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(301) & concat_CP_34_elements(302);
      gj_concat_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	296 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	551 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	294 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_sample_complete
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Sample/ack
      -- 
    ack_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_0, ack => concat_CP_34_elements(300)); -- 
    -- CP-element group 301:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	297 
    -- CP-element group 301: marked-successors 
    -- CP-element group 301: 	299 
    -- CP-element group 301:  members (8) 
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_root_address_calculated
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_offset_calculated
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_final_index_sum_regn_Update/ack
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/$entry
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/$exit
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/sum_rename_req
      -- CP-element group 301: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_876_base_plus_offset/sum_rename_ack
      -- 
    ack_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_1, ack => concat_CP_34_elements(301)); -- 
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: successors 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	299 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_sample_completed_
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/$exit
      -- CP-element group 302: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_request/ack
      -- 
    ack_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_0, ack => concat_CP_34_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	298 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	308 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	298 
    -- CP-element group 303:  members (19) 
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_update_completed_
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_877_complete/ack
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_word_addrgen/root_register_ack
      -- 
    ack_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_1, ack => concat_CP_34_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	288 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/req
      -- 
    req_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(304), ack => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0); -- 
    concat_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(306);
      gj_concat_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	310 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_update_start_
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/req
      -- 
    req_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(305), ack => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1); -- 
    concat_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(307) & concat_CP_34_elements(310);
      gj_concat_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: marked-successors 
    -- CP-element group 306: 	286 
    -- CP-element group 306: 	304 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Sample/ack
      -- 
    ack_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0, ack => concat_CP_34_elements(306)); -- 
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_881_Update/ack
      -- 
    ack_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1, ack => concat_CP_34_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	303 
    -- CP-element group 308: 	307 
    -- CP-element group 308: marked-predecessors 
    -- CP-element group 308: 	310 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/$entry
      -- CP-element group 308: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/rr
      -- 
    rr_1774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(308), ack => ptr_deref_885_load_0_req_0); -- 
    concat_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(303) & concat_CP_34_elements(307) & concat_CP_34_elements(310);
      gj_concat_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: 	337 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (5) 
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_update_start_
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/$entry
      -- CP-element group 309: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/cr
      -- 
    cr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(309), ack => ptr_deref_885_load_0_req_1); -- 
    concat_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(311) & concat_CP_34_elements(337);
      gj_concat_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310: marked-successors 
    -- CP-element group 310: 	298 
    -- CP-element group 310: 	305 
    -- CP-element group 310: 	308 
    -- CP-element group 310:  members (5) 
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/$exit
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/$exit
      -- CP-element group 310: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Sample/word_access_start/word_0/ra
      -- 
    ra_1775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_885_load_0_ack_0, ack => concat_CP_34_elements(310)); -- 
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	335 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311:  members (9) 
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/$exit
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/$exit
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/word_access_complete/word_0/ca
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/$entry
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/$exit
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/merge_req
      -- CP-element group 311: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_885_Update/ptr_deref_885_Merge/merge_ack
      -- 
    ca_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_885_load_0_ack_1, ack => concat_CP_34_elements(311)); -- 
    -- CP-element group 312:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	185 
    -- CP-element group 312: marked-predecessors 
    -- CP-element group 312: 	314 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/req
      -- 
    req_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(312), ack => W_add_outx_x1_883_delayed_1_0_887_inst_req_0); -- 
    concat_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(185) & concat_CP_34_elements(314);
      gj_concat_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: 	318 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_update_start_
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/req
      -- 
    req_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(313), ack => W_add_outx_x1_883_delayed_1_0_887_inst_req_1); -- 
    concat_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(315) & concat_CP_34_elements(318);
      gj_concat_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: successors 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	183 
    -- CP-element group 314: 	312 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Sample/ack
      -- 
    ack_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_883_delayed_1_0_887_inst_ack_0, ack => concat_CP_34_elements(314)); -- 
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	313 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_889_Update/ack
      -- 
    ack_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_883_delayed_1_0_887_inst_ack_1, ack => concat_CP_34_elements(315)); -- 
    -- CP-element group 316:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	288 
    -- CP-element group 316: 	315 
    -- CP-element group 316: marked-predecessors 
    -- CP-element group 316: 	318 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/rr
      -- 
    rr_1813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(316), ack => type_cast_893_inst_req_0); -- 
    concat_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(315) & concat_CP_34_elements(318);
      gj_concat_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: 	323 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_update_start_
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/cr
      -- 
    cr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(317), ack => type_cast_893_inst_req_1); -- 
    concat_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(319) & concat_CP_34_elements(323);
      gj_concat_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: successors 
    -- CP-element group 318: marked-successors 
    -- CP-element group 318: 	286 
    -- CP-element group 318: 	313 
    -- CP-element group 318: 	316 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Sample/ra
      -- 
    ra_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_0, ack => concat_CP_34_elements(318)); -- 
    -- CP-element group 319:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	323 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	317 
    -- CP-element group 319:  members (16) 
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/index_resize_ack
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/scale_rename_req
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scale_1/scale_rename_ack
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/req
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/index_resize_req
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resize_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_computed_1
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_scaled_1
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_893_Update/ca
      -- CP-element group 319: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_index_resized_1
      -- 
    ca_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_893_inst_ack_1, ack => concat_CP_34_elements(319)); -- 
    req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(319), ack => array_obj_ref_899_index_offset_req_0); -- 
    -- CP-element group 320:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	324 
    -- CP-element group 320: marked-predecessors 
    -- CP-element group 320: 	325 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	325 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/req
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/$entry
      -- CP-element group 320: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_sample_start_
      -- 
    req_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(320), ack => addr_of_900_final_reg_req_0); -- 
    concat_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(324) & concat_CP_34_elements(325);
      gj_concat_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	176 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	326 
    -- CP-element group 321: 	333 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	326 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/$entry
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/req
      -- CP-element group 321: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_update_start_
      -- 
    req_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(321), ack => addr_of_900_final_reg_req_1); -- 
    concat_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(326) & concat_CP_34_elements(333);
      gj_concat_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	176 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: 	325 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/req
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_update_start
      -- 
    req_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(322), ack => array_obj_ref_899_index_offset_req_1); -- 
    concat_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(324) & concat_CP_34_elements(325);
      gj_concat_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	319 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	551 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	317 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_sample_complete
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Sample/$exit
      -- 
    ack_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_899_index_offset_ack_0, ack => concat_CP_34_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	320 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (8) 
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/$entry
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/$exit
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_final_index_sum_regn_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/sum_rename_ack
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_base_plus_offset/sum_rename_req
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_root_address_calculated
      -- CP-element group 324: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_899_offset_calculated
      -- 
    ack_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_899_index_offset_ack_1, ack => concat_CP_34_elements(324)); -- 
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	320 
    -- CP-element group 325: successors 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	322 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/ack
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_request/$exit
      -- CP-element group 325: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_sample_completed_
      -- 
    ack_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_900_final_reg_ack_0, ack => concat_CP_34_elements(325)); -- 
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	321 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	331 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	321 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/ack
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_complete/$exit
      -- CP-element group 326: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_900_update_completed_
      -- 
    ack_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_900_final_reg_ack_1, ack => concat_CP_34_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	288 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	329 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_sample_start_
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/$entry
      -- CP-element group 327: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/req
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(327), ack => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0); -- 
    concat_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(329);
      gj_concat_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	330 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_update_start_
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/req
      -- CP-element group 328: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/$entry
      -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(328), ack => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1); -- 
    concat_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(330);
      gj_concat_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329: marked-successors 
    -- CP-element group 329: 	286 
    -- CP-element group 329: 	327 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Sample/ack
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0, ack => concat_CP_34_elements(329)); -- 
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	551 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	328 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/ack
      -- CP-element group 330: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_904_Update/$exit
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1, ack => concat_CP_34_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	326 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	333 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/req
      -- CP-element group 331: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_sample_start_
      -- 
    req_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(331), ack => W_arrayidx252_894_delayed_6_0_905_inst_req_0); -- 
    concat_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(326) & concat_CP_34_elements(333);
      gj_concat_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: marked-predecessors 
    -- CP-element group 332: 	334 
    -- CP-element group 332: 	337 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	334 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/req
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/$entry
      -- CP-element group 332: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_update_start_
      -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(332), ack => W_arrayidx252_894_delayed_6_0_905_inst_req_1); -- 
    concat_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(334) & concat_CP_34_elements(337);
      gj_concat_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: successors 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	321 
    -- CP-element group 333: 	331 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_sample_completed_
      -- 
    ack_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx252_894_delayed_6_0_905_inst_ack_0, ack => concat_CP_34_elements(333)); -- 
    -- CP-element group 334:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	332 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334: marked-successors 
    -- CP-element group 334: 	332 
    -- CP-element group 334:  members (19) 
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_root_address_calculated
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/sum_rename_req
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_address_calculated
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/sum_rename_ack
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/$entry
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_address_calculated
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/$entry
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/$exit
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_907_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/base_resize_req
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_addr_resize/base_resize_ack
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/$exit
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/$entry
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_plus_offset/$exit
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_base_address_resized
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/root_register_req
      -- CP-element group 334: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_word_addrgen/root_register_ack
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx252_894_delayed_6_0_905_inst_ack_1, ack => concat_CP_34_elements(334)); -- 
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	311 
    -- CP-element group 335: 	334 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	447 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (9) 
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/split_ack
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/$entry
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/$entry
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/split_req
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/$exit
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/rr
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/ptr_deref_910_Split/$entry
      -- 
    rr_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(335), ack => ptr_deref_910_store_0_req_0); -- 
    concat_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(311) & concat_CP_34_elements(334) & concat_CP_34_elements(337) & concat_CP_34_elements(447);
      gj_concat_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: marked-predecessors 
    -- CP-element group 336: 	338 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_update_start_
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/$entry
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/cr
      -- CP-element group 336: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/$entry
      -- 
    cr_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(336), ack => ptr_deref_910_store_0_req_1); -- 
    concat_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(338);
      gj_concat_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	550 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	309 
    -- CP-element group 337: 	332 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (5) 
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/ra
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/word_0/$exit
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/word_access_start/$exit
      -- CP-element group 337: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Sample/$exit
      -- 
    ra_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_910_store_0_ack_0, ack => concat_CP_34_elements(337)); -- 
    -- CP-element group 338:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	551 
    -- CP-element group 338: marked-successors 
    -- CP-element group 338: 	336 
    -- CP-element group 338:  members (5) 
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/$exit
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/ca
      -- CP-element group 338: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_Update/word_access_complete/word_0/$exit
      -- 
    ca_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_910_store_0_ack_1, ack => concat_CP_34_elements(338)); -- 
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	248 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/req
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_sample_start_
      -- 
    req_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(339), ack => W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0); -- 
    concat_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(248) & concat_CP_34_elements(341);
      gj_concat_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: marked-predecessors 
    -- CP-element group 340: 	342 
    -- CP-element group 340: 	365 
    -- CP-element group 340: 	523 
    -- CP-element group 340: 	527 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/req
      -- CP-element group 340: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_update_start_
      -- 
    req_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(340), ack => W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1); -- 
    concat_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(342) & concat_CP_34_elements(365) & concat_CP_34_elements(523) & concat_CP_34_elements(527);
      gj_concat_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	244 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_sample_completed_
      -- 
    ack_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0, ack => concat_CP_34_elements(341)); -- 
    -- CP-element group 342:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	363 
    -- CP-element group 342: 	521 
    -- CP-element group 342: 	525 
    -- CP-element group 342: marked-successors 
    -- CP-element group 342: 	340 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_915_update_completed_
      -- 
    ack_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1, ack => concat_CP_34_elements(342)); -- 
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	206 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/req
      -- CP-element group 343: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_sample_start_
      -- 
    req_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(343), ack => W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0); -- 
    concat_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(206) & concat_CP_34_elements(345);
      gj_concat_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	179 
    -- CP-element group 344: marked-predecessors 
    -- CP-element group 344: 	346 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/req
      -- CP-element group 344: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_update_start_
      -- 
    req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(344), ack => W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1); -- 
    concat_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(346);
      gj_concat_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: marked-successors 
    -- CP-element group 345: 	202 
    -- CP-element group 345: 	343 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_sample_completed_
      -- 
    ack_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0, ack => concat_CP_34_elements(345)); -- 
    -- CP-element group 346:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	551 
    -- CP-element group 346: marked-successors 
    -- CP-element group 346: 	201 
    -- CP-element group 346: 	344 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_925_update_completed_
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1, ack => concat_CP_34_elements(346)); -- 
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	185 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	349 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	349 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/req
      -- CP-element group 347: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_sample_start_
      -- 
    req_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(347), ack => W_add_outx_x1_914_delayed_1_0_933_inst_req_0); -- 
    concat_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(185) & concat_CP_34_elements(349);
      gj_concat_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	424 
    -- CP-element group 348: 	459 
    -- CP-element group 348: 	463 
    -- CP-element group 348: 	515 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/req
      -- CP-element group 348: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_update_start_
      -- 
    req_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(348), ack => W_add_outx_x1_914_delayed_1_0_933_inst_req_1); -- 
    concat_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(350) & concat_CP_34_elements(424) & concat_CP_34_elements(459) & concat_CP_34_elements(463) & concat_CP_34_elements(515);
      gj_concat_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	183 
    -- CP-element group 349: 	347 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/ack
      -- CP-element group 349: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_sample_completed_
      -- 
    ack_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_914_delayed_1_0_933_inst_ack_0, ack => concat_CP_34_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	422 
    -- CP-element group 350: 	457 
    -- CP-element group 350: 	461 
    -- CP-element group 350: 	513 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/ack
      -- CP-element group 350: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_935_update_completed_
      -- 
    ack_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_914_delayed_1_0_933_inst_ack_1, ack => concat_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	185 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	353 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/rr
      -- CP-element group 351: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_sample_start_
      -- 
    rr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(351), ack => type_cast_953_inst_req_0); -- 
    concat_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(185) & concat_CP_34_elements(353);
      gj_concat_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: marked-predecessors 
    -- CP-element group 352: 	354 
    -- CP-element group 352: 	424 
    -- CP-element group 352: 	459 
    -- CP-element group 352: 	463 
    -- CP-element group 352: 	515 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/cr
      -- CP-element group 352: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_update_start_
      -- 
    cr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(352), ack => type_cast_953_inst_req_1); -- 
    concat_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(354) & concat_CP_34_elements(424) & concat_CP_34_elements(459) & concat_CP_34_elements(463) & concat_CP_34_elements(515);
      gj_concat_cp_element_group_352 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: marked-successors 
    -- CP-element group 353: 	183 
    -- CP-element group 353: 	351 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Sample/ra
      -- CP-element group 353: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_sample_completed_
      -- 
    ra_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_0, ack => concat_CP_34_elements(353)); -- 
    -- CP-element group 354:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	422 
    -- CP-element group 354: 	457 
    -- CP-element group 354: 	461 
    -- CP-element group 354: 	513 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	352 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_953_Update/ca
      -- 
    ca_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_1, ack => concat_CP_34_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	206 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	357 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/$entry
      -- 
    rr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(355), ack => type_cast_968_inst_req_0); -- 
    concat_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(206) & concat_CP_34_elements(357);
      gj_concat_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	179 
    -- CP-element group 356: marked-predecessors 
    -- CP-element group 356: 	358 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/cr
      -- CP-element group 356: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_update_start_
      -- 
    cr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(356), ack => type_cast_968_inst_req_1); -- 
    concat_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(358);
      gj_concat_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: marked-successors 
    -- CP-element group 357: 	202 
    -- CP-element group 357: 	355 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Sample/ra
      -- CP-element group 357: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_sample_completed_
      -- 
    ra_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_0, ack => concat_CP_34_elements(357)); -- 
    -- CP-element group 358:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	551 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	201 
    -- CP-element group 358: 	356 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_968_Update/ca
      -- 
    ca_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_968_inst_ack_1, ack => concat_CP_34_elements(358)); -- 
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	248 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	361 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_sample_start_
      -- 
    rr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(359), ack => type_cast_983_inst_req_0); -- 
    concat_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(248) & concat_CP_34_elements(361);
      gj_concat_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: marked-predecessors 
    -- CP-element group 360: 	362 
    -- CP-element group 360: 	365 
    -- CP-element group 360: 	523 
    -- CP-element group 360: 	527 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/cr
      -- CP-element group 360: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_update_start_
      -- 
    cr_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(360), ack => type_cast_983_inst_req_1); -- 
    concat_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(362) & concat_CP_34_elements(365) & concat_CP_34_elements(523) & concat_CP_34_elements(527);
      gj_concat_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: marked-successors 
    -- CP-element group 361: 	244 
    -- CP-element group 361: 	359 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Sample/ra
      -- CP-element group 361: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_sample_completed_
      -- 
    ra_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_983_inst_ack_0, ack => concat_CP_34_elements(361)); -- 
    -- CP-element group 362:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362: 	521 
    -- CP-element group 362: 	525 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	360 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_Update/ca
      -- CP-element group 362: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_983_update_completed_
      -- 
    ca_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_983_inst_ack_1, ack => concat_CP_34_elements(362)); -- 
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	288 
    -- CP-element group 363: 	342 
    -- CP-element group 363: 	362 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/rr
      -- CP-element group 363: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/$entry
      -- 
    rr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(363), ack => type_cast_999_inst_req_0); -- 
    concat_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(342) & concat_CP_34_elements(362) & concat_CP_34_elements(365);
      gj_concat_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: 	385 
    -- CP-element group 364: 	389 
    -- CP-element group 364: 	393 
    -- CP-element group 364: 	397 
    -- CP-element group 364: 	503 
    -- CP-element group 364: 	519 
    -- CP-element group 364: 	531 
    -- CP-element group 364: 	543 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	366 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/cr
      -- CP-element group 364: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_update_start_
      -- 
    cr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(364), ack => type_cast_999_inst_req_1); -- 
    concat_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(385) & concat_CP_34_elements(389) & concat_CP_34_elements(393) & concat_CP_34_elements(397) & concat_CP_34_elements(503) & concat_CP_34_elements(519) & concat_CP_34_elements(531) & concat_CP_34_elements(543);
      gj_concat_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	286 
    -- CP-element group 365: 	340 
    -- CP-element group 365: 	360 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Sample/$exit
      -- 
    ra_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_0, ack => concat_CP_34_elements(365)); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	364 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	383 
    -- CP-element group 366: 	387 
    -- CP-element group 366: 	391 
    -- CP-element group 366: 	395 
    -- CP-element group 366: 	501 
    -- CP-element group 366: 	517 
    -- CP-element group 366: 	529 
    -- CP-element group 366: 	541 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/ca
      -- CP-element group 366: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_999_update_completed_
      -- 
    ca_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_1, ack => concat_CP_34_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	288 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/req
      -- CP-element group 367: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_sample_start_
      -- 
    req_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(367), ack => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0); -- 
    concat_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(369);
      gj_concat_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: marked-predecessors 
    -- CP-element group 368: 	370 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/req
      -- CP-element group 368: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_update_start_
      -- 
    req_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(368), ack => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1); -- 
    concat_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(370);
      gj_concat_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	286 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/ack
      -- CP-element group 369: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_sample_completed_
      -- 
    ack_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0, ack => concat_CP_34_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	551 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	368 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/ack
      -- CP-element group 370: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1003_update_completed_
      -- 
    ack_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1, ack => concat_CP_34_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	288 
    -- CP-element group 371: marked-predecessors 
    -- CP-element group 371: 	373 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/req
      -- 
    req_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(371), ack => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0); -- 
    concat_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(373);
      gj_concat_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: 	385 
    -- CP-element group 372: 	389 
    -- CP-element group 372: 	393 
    -- CP-element group 372: 	397 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_update_start_
      -- CP-element group 372: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/req
      -- CP-element group 372: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/$entry
      -- 
    req_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(372), ack => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1); -- 
    concat_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(374) & concat_CP_34_elements(385) & concat_CP_34_elements(389) & concat_CP_34_elements(393) & concat_CP_34_elements(397);
      gj_concat_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: successors 
    -- CP-element group 373: marked-successors 
    -- CP-element group 373: 	286 
    -- CP-element group 373: 	371 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_sample_completed_
      -- CP-element group 373: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/ack
      -- CP-element group 373: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Sample/$exit
      -- 
    ack_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0, ack => concat_CP_34_elements(373)); -- 
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	383 
    -- CP-element group 374: 	387 
    -- CP-element group 374: 	391 
    -- CP-element group 374: 	395 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_update_completed_
      -- CP-element group 374: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/ack
      -- CP-element group 374: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1012_Update/$exit
      -- 
    ack_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1, ack => concat_CP_34_elements(374)); -- 
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	288 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/req
      -- CP-element group 375: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_sample_start_
      -- 
    req_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(375), ack => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0); -- 
    concat_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(377);
      gj_concat_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: 	503 
    -- CP-element group 376: 	519 
    -- CP-element group 376: 	531 
    -- CP-element group 376: 	543 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_update_start_
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/req
      -- 
    req_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(376), ack => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1); -- 
    concat_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_CP_34_elements(378) & concat_CP_34_elements(503) & concat_CP_34_elements(519) & concat_CP_34_elements(531) & concat_CP_34_elements(543);
      gj_concat_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	286 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Sample/ack
      -- CP-element group 377: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_sample_completed_
      -- 
    ack_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0, ack => concat_CP_34_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	501 
    -- CP-element group 378: 	517 
    -- CP-element group 378: 	529 
    -- CP-element group 378: 	541 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1020_Update/ack
      -- 
    ack_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1, ack => concat_CP_34_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	269 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/req
      -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(379), ack => W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0); -- 
    concat_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(269) & concat_CP_34_elements(381);
      gj_concat_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: 	385 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_update_start_
      -- CP-element group 380: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/req
      -- CP-element group 380: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/$entry
      -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(380), ack => W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1); -- 
    concat_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(382) & concat_CP_34_elements(385);
      gj_concat_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	265 
    -- CP-element group 381: 	379 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Sample/ack
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0, ack => concat_CP_34_elements(381)); -- 
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/ack
      -- CP-element group 382: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1032_Update/$exit
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1, ack => concat_CP_34_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	366 
    -- CP-element group 383: 	374 
    -- CP-element group 383: 	382 
    -- CP-element group 383: marked-predecessors 
    -- CP-element group 383: 	385 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	385 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/rr
      -- CP-element group 383: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_sample_start_
      -- 
    rr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(383), ack => type_cast_1036_inst_req_0); -- 
    concat_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(374) & concat_CP_34_elements(382) & concat_CP_34_elements(385);
      gj_concat_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: 	405 
    -- CP-element group 384: 	416 
    -- CP-element group 384: 	428 
    -- CP-element group 384: 	439 
    -- CP-element group 384: 	475 
    -- CP-element group 384: 	479 
    -- CP-element group 384: 	483 
    -- CP-element group 384: 	487 
    -- CP-element group 384: 	491 
    -- CP-element group 384: 	495 
    -- CP-element group 384: 	507 
    -- CP-element group 384: 	511 
    -- CP-element group 384: 	535 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_update_start_
      -- 
    cr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(384), ack => type_cast_1036_inst_req_1); -- 
    concat_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(405) & concat_CP_34_elements(416) & concat_CP_34_elements(428) & concat_CP_34_elements(439) & concat_CP_34_elements(475) & concat_CP_34_elements(479) & concat_CP_34_elements(483) & concat_CP_34_elements(487) & concat_CP_34_elements(491) & concat_CP_34_elements(495) & concat_CP_34_elements(507) & concat_CP_34_elements(511) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	383 
    -- CP-element group 385: successors 
    -- CP-element group 385: marked-successors 
    -- CP-element group 385: 	364 
    -- CP-element group 385: 	372 
    -- CP-element group 385: 	380 
    -- CP-element group 385: 	383 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/ra
      -- CP-element group 385: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_sample_completed_
      -- 
    ra_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_0, ack => concat_CP_34_elements(385)); -- 
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	403 
    -- CP-element group 386: 	414 
    -- CP-element group 386: 	426 
    -- CP-element group 386: 	437 
    -- CP-element group 386: 	473 
    -- CP-element group 386: 	477 
    -- CP-element group 386: 	481 
    -- CP-element group 386: 	485 
    -- CP-element group 386: 	489 
    -- CP-element group 386: 	493 
    -- CP-element group 386: 	505 
    -- CP-element group 386: 	509 
    -- CP-element group 386: 	533 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/ca
      -- CP-element group 386: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1036_update_completed_
      -- 
    ca_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1036_inst_ack_1, ack => concat_CP_34_elements(386)); -- 
    -- CP-element group 387:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	366 
    -- CP-element group 387: 	374 
    -- CP-element group 387: marked-predecessors 
    -- CP-element group 387: 	389 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	389 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/req
      -- CP-element group 387: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/$entry
      -- 
    req_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(387), ack => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0); -- 
    concat_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(374) & concat_CP_34_elements(389);
      gj_concat_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: marked-predecessors 
    -- CP-element group 388: 	390 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	390 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_update_start_
      -- CP-element group 388: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/req
      -- CP-element group 388: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/$entry
      -- 
    req_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(388), ack => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1); -- 
    concat_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(390);
      gj_concat_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	387 
    -- CP-element group 389: successors 
    -- CP-element group 389: marked-successors 
    -- CP-element group 389: 	364 
    -- CP-element group 389: 	372 
    -- CP-element group 389: 	387 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/ack
      -- CP-element group 389: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Sample/$exit
      -- 
    ack_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0, ack => concat_CP_34_elements(389)); -- 
    -- CP-element group 390:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	388 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	551 
    -- CP-element group 390: marked-successors 
    -- CP-element group 390: 	388 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/ack
      -- CP-element group 390: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1040_update_completed_
      -- 
    ack_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1, ack => concat_CP_34_elements(390)); -- 
    -- CP-element group 391:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	366 
    -- CP-element group 391: 	374 
    -- CP-element group 391: marked-predecessors 
    -- CP-element group 391: 	393 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	393 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/req
      -- CP-element group 391: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/$entry
      -- 
    req_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(391), ack => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0); -- 
    concat_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(374) & concat_CP_34_elements(393);
      gj_concat_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: marked-predecessors 
    -- CP-element group 392: 	394 
    -- CP-element group 392: 	405 
    -- CP-element group 392: 	416 
    -- CP-element group 392: 	428 
    -- CP-element group 392: 	439 
    -- CP-element group 392: 	475 
    -- CP-element group 392: 	479 
    -- CP-element group 392: 	483 
    -- CP-element group 392: 	487 
    -- CP-element group 392: 	491 
    -- CP-element group 392: 	495 
    -- CP-element group 392: 	507 
    -- CP-element group 392: 	511 
    -- CP-element group 392: 	535 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	394 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_update_start_
      -- CP-element group 392: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/req
      -- CP-element group 392: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/$entry
      -- 
    req_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(392), ack => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1); -- 
    concat_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= concat_CP_34_elements(394) & concat_CP_34_elements(405) & concat_CP_34_elements(416) & concat_CP_34_elements(428) & concat_CP_34_elements(439) & concat_CP_34_elements(475) & concat_CP_34_elements(479) & concat_CP_34_elements(483) & concat_CP_34_elements(487) & concat_CP_34_elements(491) & concat_CP_34_elements(495) & concat_CP_34_elements(507) & concat_CP_34_elements(511) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_392 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	391 
    -- CP-element group 393: successors 
    -- CP-element group 393: marked-successors 
    -- CP-element group 393: 	364 
    -- CP-element group 393: 	372 
    -- CP-element group 393: 	391 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/ack
      -- CP-element group 393: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Sample/$exit
      -- 
    ack_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0, ack => concat_CP_34_elements(393)); -- 
    -- CP-element group 394:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	392 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	403 
    -- CP-element group 394: 	414 
    -- CP-element group 394: 	426 
    -- CP-element group 394: 	437 
    -- CP-element group 394: 	473 
    -- CP-element group 394: 	477 
    -- CP-element group 394: 	481 
    -- CP-element group 394: 	485 
    -- CP-element group 394: 	489 
    -- CP-element group 394: 	493 
    -- CP-element group 394: 	505 
    -- CP-element group 394: 	509 
    -- CP-element group 394: 	533 
    -- CP-element group 394: marked-successors 
    -- CP-element group 394: 	392 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/ack
      -- CP-element group 394: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1049_Update/$exit
      -- 
    ack_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1, ack => concat_CP_34_elements(394)); -- 
    -- CP-element group 395:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	366 
    -- CP-element group 395: 	374 
    -- CP-element group 395: marked-predecessors 
    -- CP-element group 395: 	397 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/req
      -- CP-element group 395: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/$entry
      -- 
    req_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(395), ack => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0); -- 
    concat_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(374) & concat_CP_34_elements(397);
      gj_concat_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: marked-predecessors 
    -- CP-element group 396: 	398 
    -- CP-element group 396: 	475 
    -- CP-element group 396: 	479 
    -- CP-element group 396: 	483 
    -- CP-element group 396: 	487 
    -- CP-element group 396: 	491 
    -- CP-element group 396: 	495 
    -- CP-element group 396: 	507 
    -- CP-element group 396: 	511 
    -- CP-element group 396: 	535 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	398 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_update_start_
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/req
      -- 
    req_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(396), ack => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1); -- 
    concat_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= concat_CP_34_elements(398) & concat_CP_34_elements(475) & concat_CP_34_elements(479) & concat_CP_34_elements(483) & concat_CP_34_elements(487) & concat_CP_34_elements(491) & concat_CP_34_elements(495) & concat_CP_34_elements(507) & concat_CP_34_elements(511) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397: marked-successors 
    -- CP-element group 397: 	364 
    -- CP-element group 397: 	372 
    -- CP-element group 397: 	395 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/ack
      -- CP-element group 397: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Sample/$exit
      -- 
    ack_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0, ack => concat_CP_34_elements(397)); -- 
    -- CP-element group 398:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	473 
    -- CP-element group 398: 	477 
    -- CP-element group 398: 	481 
    -- CP-element group 398: 	485 
    -- CP-element group 398: 	489 
    -- CP-element group 398: 	493 
    -- CP-element group 398: 	505 
    -- CP-element group 398: 	509 
    -- CP-element group 398: 	533 
    -- CP-element group 398: marked-successors 
    -- CP-element group 398: 	396 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_Update/ack
      -- CP-element group 398: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1057_update_completed_
      -- 
    ack_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1, ack => concat_CP_34_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	227 
    -- CP-element group 399: marked-predecessors 
    -- CP-element group 399: 	401 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	401 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_sample_start_
      -- 
    req_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(399), ack => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0); -- 
    concat_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(227) & concat_CP_34_elements(401);
      gj_concat_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: marked-predecessors 
    -- CP-element group 400: 	402 
    -- CP-element group 400: 	405 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_update_start_
      -- CP-element group 400: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/req
      -- 
    req_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(400), ack => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1); -- 
    concat_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(402) & concat_CP_34_elements(405);
      gj_concat_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	399 
    -- CP-element group 401: successors 
    -- CP-element group 401: marked-successors 
    -- CP-element group 401: 	223 
    -- CP-element group 401: 	399 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/ack
      -- CP-element group 401: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_sample_completed_
      -- 
    ack_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0, ack => concat_CP_34_elements(401)); -- 
    -- CP-element group 402:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402: marked-successors 
    -- CP-element group 402: 	400 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1069_Update/ack
      -- 
    ack_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1, ack => concat_CP_34_elements(402)); -- 
    -- CP-element group 403:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	386 
    -- CP-element group 403: 	394 
    -- CP-element group 403: 	402 
    -- CP-element group 403: marked-predecessors 
    -- CP-element group 403: 	405 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/$entry
      -- 
    rr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(403), ack => type_cast_1073_inst_req_0); -- 
    concat_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(402) & concat_CP_34_elements(405);
      gj_concat_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: marked-predecessors 
    -- CP-element group 404: 	406 
    -- CP-element group 404: 	410 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	406 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_update_start_
      -- 
    cr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(404), ack => type_cast_1073_inst_req_1); -- 
    concat_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(406) & concat_CP_34_elements(410);
      gj_concat_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: successors 
    -- CP-element group 405: marked-successors 
    -- CP-element group 405: 	384 
    -- CP-element group 405: 	392 
    -- CP-element group 405: 	400 
    -- CP-element group 405: 	403 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Sample/ra
      -- 
    ra_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_0, ack => concat_CP_34_elements(405)); -- 
    -- CP-element group 406:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	404 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	410 
    -- CP-element group 406: marked-successors 
    -- CP-element group 406: 	404 
    -- CP-element group 406:  members (16) 
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_update_completed_
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1073_Update/ca
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resized_1
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scaled_1
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_computed_1
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/$entry
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/$exit
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/index_resize_req
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_resize_1/index_resize_ack
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/$entry
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/$exit
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/scale_rename_req
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_index_scale_1/scale_rename_ack
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/req
      -- 
    ca_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_1, ack => concat_CP_34_elements(406)); -- 
    req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(406), ack => array_obj_ref_1079_index_offset_req_0); -- 
    -- CP-element group 407:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	411 
    -- CP-element group 407: marked-predecessors 
    -- CP-element group 407: 	412 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	412 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/$entry
      -- CP-element group 407: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/req
      -- 
    req_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(407), ack => addr_of_1080_final_reg_req_0); -- 
    concat_cp_element_group_407: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_407"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(411) & concat_CP_34_elements(412);
      gj_concat_cp_element_group_407 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(407), clk => clk, reset => reset); --
    end block;
    -- CP-element group 408:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	176 
    -- CP-element group 408: marked-predecessors 
    -- CP-element group 408: 	413 
    -- CP-element group 408: 	420 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	413 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_update_start_
      -- CP-element group 408: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/$entry
      -- CP-element group 408: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/req
      -- 
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(408), ack => addr_of_1080_final_reg_req_1); -- 
    concat_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(413) & concat_CP_34_elements(420);
      gj_concat_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	176 
    -- CP-element group 409: marked-predecessors 
    -- CP-element group 409: 	411 
    -- CP-element group 409: 	412 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_update_start
      -- CP-element group 409: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/req
      -- 
    req_2211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(409), ack => array_obj_ref_1079_index_offset_req_1); -- 
    concat_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(411) & concat_CP_34_elements(412);
      gj_concat_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	406 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	551 
    -- CP-element group 410: marked-successors 
    -- CP-element group 410: 	404 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_sample_complete
      -- CP-element group 410: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Sample/ack
      -- 
    ack_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_0, ack => concat_CP_34_elements(410)); -- 
    -- CP-element group 411:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	409 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	407 
    -- CP-element group 411: marked-successors 
    -- CP-element group 411: 	409 
    -- CP-element group 411:  members (8) 
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_root_address_calculated
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_offset_calculated
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_final_index_sum_regn_Update/ack
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/$entry
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/$exit
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_req
      -- CP-element group 411: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_ack
      -- 
    ack_2212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_1, ack => concat_CP_34_elements(411)); -- 
    -- CP-element group 412:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	407 
    -- CP-element group 412: successors 
    -- CP-element group 412: marked-successors 
    -- CP-element group 412: 	407 
    -- CP-element group 412: 	409 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/$exit
      -- CP-element group 412: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_request/ack
      -- 
    ack_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_0, ack => concat_CP_34_elements(412)); -- 
    -- CP-element group 413:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	408 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	418 
    -- CP-element group 413: marked-successors 
    -- CP-element group 413: 	408 
    -- CP-element group 413:  members (19) 
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/$exit
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1080_complete/ack
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_address_calculated
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_address_calculated
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_root_address_calculated
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_address_resized
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/$entry
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/$exit
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/base_resize_req
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_addr_resize/base_resize_ack
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/$entry
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/$exit
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/sum_rename_req
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_base_plus_offset/sum_rename_ack
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/$entry
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/$exit
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/root_register_req
      -- CP-element group 413: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_word_addrgen/root_register_ack
      -- 
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_1, ack => concat_CP_34_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	386 
    -- CP-element group 414: 	394 
    -- CP-element group 414: marked-predecessors 
    -- CP-element group 414: 	416 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	416 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_sample_start_
      -- CP-element group 414: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/req
      -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(414), ack => W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_0); -- 
    concat_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(416);
      gj_concat_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: marked-predecessors 
    -- CP-element group 415: 	417 
    -- CP-element group 415: 	420 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	417 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_update_start_
      -- CP-element group 415: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/req
      -- 
    req_2240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(415), ack => W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_1); -- 
    concat_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(417) & concat_CP_34_elements(420);
      gj_concat_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416: marked-successors 
    -- CP-element group 416: 	384 
    -- CP-element group 416: 	392 
    -- CP-element group 416: 	414 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Sample/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_0, ack => concat_CP_34_elements(416)); -- 
    -- CP-element group 417:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	415 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417: marked-successors 
    -- CP-element group 417: 	415 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1084_Update/ack
      -- 
    ack_2241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_1, ack => concat_CP_34_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	413 
    -- CP-element group 418: 	417 
    -- CP-element group 418: marked-predecessors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/$entry
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/$entry
      -- CP-element group 418: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/rr
      -- 
    rr_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(418), ack => ptr_deref_1088_load_0_req_0); -- 
    concat_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(413) & concat_CP_34_elements(417) & concat_CP_34_elements(420);
      gj_concat_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: marked-predecessors 
    -- CP-element group 419: 	421 
    -- CP-element group 419: 	447 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	421 
    -- CP-element group 419:  members (5) 
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_update_start_
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/$entry
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/$entry
      -- CP-element group 419: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/cr
      -- 
    cr_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(419), ack => ptr_deref_1088_load_0_req_1); -- 
    concat_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(421) & concat_CP_34_elements(447);
      gj_concat_cp_element_group_419 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420: marked-successors 
    -- CP-element group 420: 	408 
    -- CP-element group 420: 	415 
    -- CP-element group 420: 	418 
    -- CP-element group 420:  members (5) 
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/$exit
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/$exit
      -- CP-element group 420: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Sample/word_access_start/word_0/ra
      -- 
    ra_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_load_0_ack_0, ack => concat_CP_34_elements(420)); -- 
    -- CP-element group 421:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	419 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	445 
    -- CP-element group 421: marked-successors 
    -- CP-element group 421: 	419 
    -- CP-element group 421:  members (9) 
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/$exit
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/$exit
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/word_access_complete/word_0/ca
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/$entry
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/$exit
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/merge_req
      -- CP-element group 421: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1088_Update/ptr_deref_1088_Merge/merge_ack
      -- 
    ca_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_load_0_ack_1, ack => concat_CP_34_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	288 
    -- CP-element group 422: 	350 
    -- CP-element group 422: 	354 
    -- CP-element group 422: marked-predecessors 
    -- CP-element group 422: 	424 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/$entry
      -- CP-element group 422: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/req
      -- 
    req_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(422), ack => W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0); -- 
    concat_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(350) & concat_CP_34_elements(354) & concat_CP_34_elements(424);
      gj_concat_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: marked-predecessors 
    -- CP-element group 423: 	425 
    -- CP-element group 423: 	428 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	425 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_update_start_
      -- CP-element group 423: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/req
      -- 
    req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(423), ack => W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1); -- 
    concat_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(425) & concat_CP_34_elements(428);
      gj_concat_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: successors 
    -- CP-element group 424: marked-successors 
    -- CP-element group 424: 	286 
    -- CP-element group 424: 	348 
    -- CP-element group 424: 	352 
    -- CP-element group 424: 	422 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Sample/ack
      -- 
    ack_2300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0, ack => concat_CP_34_elements(424)); -- 
    -- CP-element group 425:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	423 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425: marked-successors 
    -- CP-element group 425: 	423 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1092_Update/ack
      -- 
    ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1, ack => concat_CP_34_elements(425)); -- 
    -- CP-element group 426:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	386 
    -- CP-element group 426: 	394 
    -- CP-element group 426: 	425 
    -- CP-element group 426: marked-predecessors 
    -- CP-element group 426: 	428 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/rr
      -- 
    rr_2313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(426), ack => type_cast_1096_inst_req_0); -- 
    concat_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(425) & concat_CP_34_elements(428);
      gj_concat_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: marked-predecessors 
    -- CP-element group 427: 	429 
    -- CP-element group 427: 	433 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_update_start_
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/cr
      -- 
    cr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(427), ack => type_cast_1096_inst_req_1); -- 
    concat_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(429) & concat_CP_34_elements(433);
      gj_concat_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: marked-successors 
    -- CP-element group 428: 	384 
    -- CP-element group 428: 	392 
    -- CP-element group 428: 	423 
    -- CP-element group 428: 	426 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Sample/ra
      -- 
    ra_2314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_0, ack => concat_CP_34_elements(428)); -- 
    -- CP-element group 429:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	433 
    -- CP-element group 429: marked-successors 
    -- CP-element group 429: 	427 
    -- CP-element group 429:  members (16) 
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1096_Update/ca
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resized_1
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scaled_1
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_computed_1
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/$entry
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/$exit
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/index_resize_req
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_resize_1/index_resize_ack
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/$entry
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/$exit
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/scale_rename_req
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_index_scale_1/scale_rename_ack
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/req
      -- 
    ca_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1096_inst_ack_1, ack => concat_CP_34_elements(429)); -- 
    req_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(429), ack => array_obj_ref_1102_index_offset_req_0); -- 
    -- CP-element group 430:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	434 
    -- CP-element group 430: marked-predecessors 
    -- CP-element group 430: 	435 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	435 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/$entry
      -- CP-element group 430: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/req
      -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(430), ack => addr_of_1103_final_reg_req_0); -- 
    concat_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(434) & concat_CP_34_elements(435);
      gj_concat_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	176 
    -- CP-element group 431: marked-predecessors 
    -- CP-element group 431: 	436 
    -- CP-element group 431: 	443 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	436 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_update_start_
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/$entry
      -- CP-element group 431: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/req
      -- 
    req_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(431), ack => addr_of_1103_final_reg_req_1); -- 
    concat_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(436) & concat_CP_34_elements(443);
      gj_concat_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	176 
    -- CP-element group 432: marked-predecessors 
    -- CP-element group 432: 	434 
    -- CP-element group 432: 	435 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	434 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_update_start
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/req
      -- 
    req_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(432), ack => array_obj_ref_1102_index_offset_req_1); -- 
    concat_cp_element_group_432: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_432"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(176) & concat_CP_34_elements(434) & concat_CP_34_elements(435);
      gj_concat_cp_element_group_432 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(432), clk => clk, reset => reset); --
    end block;
    -- CP-element group 433:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	429 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	551 
    -- CP-element group 433: marked-successors 
    -- CP-element group 433: 	427 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_sample_complete
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Sample/ack
      -- 
    ack_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1102_index_offset_ack_0, ack => concat_CP_34_elements(433)); -- 
    -- CP-element group 434:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	432 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	430 
    -- CP-element group 434: marked-successors 
    -- CP-element group 434: 	432 
    -- CP-element group 434:  members (8) 
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_root_address_calculated
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_offset_calculated
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_final_index_sum_regn_Update/ack
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/$entry
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/$exit
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/sum_rename_req
      -- CP-element group 434: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/array_obj_ref_1102_base_plus_offset/sum_rename_ack
      -- 
    ack_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1102_index_offset_ack_1, ack => concat_CP_34_elements(434)); -- 
    -- CP-element group 435:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	430 
    -- CP-element group 435: successors 
    -- CP-element group 435: marked-successors 
    -- CP-element group 435: 	430 
    -- CP-element group 435: 	432 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/$exit
      -- CP-element group 435: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_request/ack
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1103_final_reg_ack_0, ack => concat_CP_34_elements(435)); -- 
    -- CP-element group 436:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	431 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	441 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	431 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/$exit
      -- CP-element group 436: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/addr_of_1103_complete/ack
      -- 
    ack_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1103_final_reg_ack_1, ack => concat_CP_34_elements(436)); -- 
    -- CP-element group 437:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	386 
    -- CP-element group 437: 	394 
    -- CP-element group 437: marked-predecessors 
    -- CP-element group 437: 	439 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	439 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/req
      -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(437), ack => W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_0); -- 
    concat_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(439);
      gj_concat_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	440 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	440 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_update_start_
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/req
      -- 
    req_2378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(438), ack => W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_1); -- 
    concat_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(440);
      gj_concat_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	437 
    -- CP-element group 439: successors 
    -- CP-element group 439: marked-successors 
    -- CP-element group 439: 	384 
    -- CP-element group 439: 	392 
    -- CP-element group 439: 	437 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Sample/ack
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_0, ack => concat_CP_34_elements(439)); -- 
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	551 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	438 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1107_Update/ack
      -- 
    ack_2379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_1, ack => concat_CP_34_elements(440)); -- 
    -- CP-element group 441:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	436 
    -- CP-element group 441: marked-predecessors 
    -- CP-element group 441: 	443 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	443 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_sample_start_
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/$entry
      -- CP-element group 441: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/req
      -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(441), ack => W_arrayidx278_1043_delayed_6_0_1108_inst_req_0); -- 
    concat_cp_element_group_441: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_441"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(436) & concat_CP_34_elements(443);
      gj_concat_cp_element_group_441 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(441), clk => clk, reset => reset); --
    end block;
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	444 
    -- CP-element group 442: 	447 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_update_start_
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/req
      -- 
    req_2392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(442), ack => W_arrayidx278_1043_delayed_6_0_1108_inst_req_1); -- 
    concat_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(444) & concat_CP_34_elements(447);
      gj_concat_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	441 
    -- CP-element group 443: successors 
    -- CP-element group 443: marked-successors 
    -- CP-element group 443: 	431 
    -- CP-element group 443: 	441 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_sample_completed_
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Sample/ack
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx278_1043_delayed_6_0_1108_inst_ack_0, ack => concat_CP_34_elements(443)); -- 
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	442 
    -- CP-element group 444:  members (19) 
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_update_completed_
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1110_Update/ack
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_address_calculated
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_address_calculated
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_root_address_calculated
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_address_resized
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/$entry
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/$exit
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/base_resize_req
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_addr_resize/base_resize_ack
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/$entry
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/$exit
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/sum_rename_req
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_base_plus_offset/sum_rename_ack
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/$entry
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/$exit
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/root_register_req
      -- CP-element group 444: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_word_addrgen/root_register_ack
      -- 
    ack_2393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx278_1043_delayed_6_0_1108_inst_ack_1, ack => concat_CP_34_elements(444)); -- 
    -- CP-element group 445:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	421 
    -- CP-element group 445: 	444 
    -- CP-element group 445: 	550 
    -- CP-element group 445: marked-predecessors 
    -- CP-element group 445: 	447 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	447 
    -- CP-element group 445:  members (9) 
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/$exit
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/split_req
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/ptr_deref_1113_Split/split_ack
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/$entry
      -- CP-element group 445: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/rr
      -- 
    rr_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(445), ack => ptr_deref_1113_store_0_req_0); -- 
    concat_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(421) & concat_CP_34_elements(444) & concat_CP_34_elements(550) & concat_CP_34_elements(447);
      gj_concat_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: marked-predecessors 
    -- CP-element group 446: 	448 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (5) 
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_update_start_
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/$entry
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/$entry
      -- CP-element group 446: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/cr
      -- 
    cr_2442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(446), ack => ptr_deref_1113_store_0_req_1); -- 
    concat_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(448);
      gj_concat_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	445 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	551 
    -- CP-element group 447: marked-successors 
    -- CP-element group 447: 	335 
    -- CP-element group 447: 	419 
    -- CP-element group 447: 	442 
    -- CP-element group 447: 	445 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ring_reenable_memory_space_2
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/$exit
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/$exit
      -- CP-element group 447: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Sample/word_access_start/word_0/ra
      -- 
    ra_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_store_0_ack_0, ack => concat_CP_34_elements(447)); -- 
    -- CP-element group 448:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	551 
    -- CP-element group 448: marked-successors 
    -- CP-element group 448: 	446 
    -- CP-element group 448:  members (5) 
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/$exit
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/$exit
      -- CP-element group 448: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_1113_Update/word_access_complete/word_0/ca
      -- 
    ca_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_store_0_ack_1, ack => concat_CP_34_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	269 
    -- CP-element group 449: marked-predecessors 
    -- CP-element group 449: 	451 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	451 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/req
      -- 
    req_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(449), ack => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0); -- 
    concat_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(269) & concat_CP_34_elements(451);
      gj_concat_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: marked-predecessors 
    -- CP-element group 450: 	452 
    -- CP-element group 450: 	475 
    -- CP-element group 450: 	535 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	452 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_update_start_
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/req
      -- 
    req_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(450), ack => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1); -- 
    concat_cp_element_group_450: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_450"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(452) & concat_CP_34_elements(475) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_450 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(450), clk => clk, reset => reset); --
    end block;
    -- CP-element group 451:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: marked-successors 
    -- CP-element group 451: 	265 
    -- CP-element group 451: 	449 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_sample_completed_
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Sample/ack
      -- 
    ack_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0, ack => concat_CP_34_elements(451)); -- 
    -- CP-element group 452:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	473 
    -- CP-element group 452: 	533 
    -- CP-element group 452: marked-successors 
    -- CP-element group 452: 	450 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_update_completed_
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1118_Update/ack
      -- 
    ack_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1, ack => concat_CP_34_elements(452)); -- 
    -- CP-element group 453:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	227 
    -- CP-element group 453: marked-predecessors 
    -- CP-element group 453: 	455 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	455 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_sample_start_
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/$entry
      -- CP-element group 453: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/req
      -- 
    req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(453), ack => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0); -- 
    concat_cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_453"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(227) & concat_CP_34_elements(455);
      gj_concat_cp_element_group_453 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 454:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: marked-predecessors 
    -- CP-element group 454: 	456 
    -- CP-element group 454: 	491 
    -- CP-element group 454: 	495 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_update_start_
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/req
      -- 
    req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(454), ack => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1); -- 
    concat_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(456) & concat_CP_34_elements(491) & concat_CP_34_elements(495);
      gj_concat_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: successors 
    -- CP-element group 455: marked-successors 
    -- CP-element group 455: 	223 
    -- CP-element group 455: 	453 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Sample/ack
      -- 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0, ack => concat_CP_34_elements(455)); -- 
    -- CP-element group 456:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	489 
    -- CP-element group 456: 	493 
    -- CP-element group 456: marked-successors 
    -- CP-element group 456: 	454 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1128_Update/ack
      -- 
    ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1, ack => concat_CP_34_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	288 
    -- CP-element group 457: 	350 
    -- CP-element group 457: 	354 
    -- CP-element group 457: marked-predecessors 
    -- CP-element group 457: 	459 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	459 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/req
      -- 
    req_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(457), ack => W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0); -- 
    concat_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(350) & concat_CP_34_elements(354) & concat_CP_34_elements(459);
      gj_concat_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: marked-predecessors 
    -- CP-element group 458: 	460 
    -- CP-element group 458: 	507 
    -- CP-element group 458: 	511 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	460 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_update_start_
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/req
      -- 
    req_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(458), ack => W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1); -- 
    concat_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(460) & concat_CP_34_elements(507) & concat_CP_34_elements(511);
      gj_concat_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: successors 
    -- CP-element group 459: marked-successors 
    -- CP-element group 459: 	286 
    -- CP-element group 459: 	348 
    -- CP-element group 459: 	352 
    -- CP-element group 459: 	457 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Sample/ack
      -- 
    ack_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0, ack => concat_CP_34_elements(459)); -- 
    -- CP-element group 460:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	505 
    -- CP-element group 460: 	509 
    -- CP-element group 460: marked-successors 
    -- CP-element group 460: 	458 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1138_Update/ack
      -- 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1, ack => concat_CP_34_elements(460)); -- 
    -- CP-element group 461:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	288 
    -- CP-element group 461: 	350 
    -- CP-element group 461: 	354 
    -- CP-element group 461: marked-predecessors 
    -- CP-element group 461: 	463 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	463 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/rr
      -- 
    rr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(461), ack => type_cast_1156_inst_req_0); -- 
    concat_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(350) & concat_CP_34_elements(354) & concat_CP_34_elements(463);
      gj_concat_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: marked-predecessors 
    -- CP-element group 462: 	464 
    -- CP-element group 462: 	507 
    -- CP-element group 462: 	511 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_update_start_
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/cr
      -- 
    cr_2498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(462), ack => type_cast_1156_inst_req_1); -- 
    concat_cp_element_group_462: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_462"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(464) & concat_CP_34_elements(507) & concat_CP_34_elements(511);
      gj_concat_cp_element_group_462 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 463:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	461 
    -- CP-element group 463: successors 
    -- CP-element group 463: marked-successors 
    -- CP-element group 463: 	286 
    -- CP-element group 463: 	348 
    -- CP-element group 463: 	352 
    -- CP-element group 463: 	461 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_sample_completed_
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Sample/ra
      -- 
    ra_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_0, ack => concat_CP_34_elements(463)); -- 
    -- CP-element group 464:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	505 
    -- CP-element group 464: 	509 
    -- CP-element group 464: marked-successors 
    -- CP-element group 464: 	462 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_update_completed_
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1156_Update/ca
      -- 
    ca_2499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1156_inst_ack_1, ack => concat_CP_34_elements(464)); -- 
    -- CP-element group 465:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	227 
    -- CP-element group 465: marked-predecessors 
    -- CP-element group 465: 	467 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	467 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/rr
      -- 
    rr_2507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(465), ack => type_cast_1171_inst_req_0); -- 
    concat_cp_element_group_465: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_465"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(227) & concat_CP_34_elements(467);
      gj_concat_cp_element_group_465 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(465), clk => clk, reset => reset); --
    end block;
    -- CP-element group 466:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: marked-predecessors 
    -- CP-element group 466: 	468 
    -- CP-element group 466: 	491 
    -- CP-element group 466: 	495 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_update_start_
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/$entry
      -- CP-element group 466: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/cr
      -- 
    cr_2512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(466), ack => type_cast_1171_inst_req_1); -- 
    concat_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(468) & concat_CP_34_elements(491) & concat_CP_34_elements(495);
      gj_concat_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	465 
    -- CP-element group 467: successors 
    -- CP-element group 467: marked-successors 
    -- CP-element group 467: 	223 
    -- CP-element group 467: 	465 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Sample/ra
      -- 
    ra_2508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => concat_CP_34_elements(467)); -- 
    -- CP-element group 468:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	489 
    -- CP-element group 468: 	493 
    -- CP-element group 468: marked-successors 
    -- CP-element group 468: 	466 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1171_Update/ca
      -- 
    ca_2513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => concat_CP_34_elements(468)); -- 
    -- CP-element group 469:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	269 
    -- CP-element group 469: marked-predecessors 
    -- CP-element group 469: 	471 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	471 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/rr
      -- 
    rr_2521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(469), ack => type_cast_1186_inst_req_0); -- 
    concat_cp_element_group_469: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_469"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(269) & concat_CP_34_elements(471);
      gj_concat_cp_element_group_469 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(469), clk => clk, reset => reset); --
    end block;
    -- CP-element group 470:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: marked-predecessors 
    -- CP-element group 470: 	472 
    -- CP-element group 470: 	475 
    -- CP-element group 470: 	535 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	472 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_update_start_
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/$entry
      -- CP-element group 470: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/cr
      -- 
    cr_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(470), ack => type_cast_1186_inst_req_1); -- 
    concat_cp_element_group_470: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_470"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(472) & concat_CP_34_elements(475) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_470 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(470), clk => clk, reset => reset); --
    end block;
    -- CP-element group 471:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	469 
    -- CP-element group 471: successors 
    -- CP-element group 471: marked-successors 
    -- CP-element group 471: 	265 
    -- CP-element group 471: 	469 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_sample_completed_
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Sample/ra
      -- 
    ra_2522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_0, ack => concat_CP_34_elements(471)); -- 
    -- CP-element group 472:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	470 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472: 	533 
    -- CP-element group 472: marked-successors 
    -- CP-element group 472: 	470 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_update_completed_
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1186_Update/ca
      -- 
    ca_2527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_1, ack => concat_CP_34_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	386 
    -- CP-element group 473: 	394 
    -- CP-element group 473: 	398 
    -- CP-element group 473: 	452 
    -- CP-element group 473: 	472 
    -- CP-element group 473: marked-predecessors 
    -- CP-element group 473: 	475 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	475 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_sample_start_
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/$entry
      -- CP-element group 473: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/rr
      -- 
    rr_2535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(473), ack => type_cast_1202_inst_req_0); -- 
    concat_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(452) & concat_CP_34_elements(472) & concat_CP_34_elements(475);
      gj_concat_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	179 
    -- CP-element group 474: marked-predecessors 
    -- CP-element group 474: 	476 
    -- CP-element group 474: 	547 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	476 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_update_start_
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/$entry
      -- CP-element group 474: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/cr
      -- 
    cr_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(474), ack => type_cast_1202_inst_req_1); -- 
    concat_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(476) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	473 
    -- CP-element group 475: successors 
    -- CP-element group 475: marked-successors 
    -- CP-element group 475: 	384 
    -- CP-element group 475: 	392 
    -- CP-element group 475: 	396 
    -- CP-element group 475: 	450 
    -- CP-element group 475: 	470 
    -- CP-element group 475: 	473 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_sample_completed_
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/$exit
      -- CP-element group 475: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Sample/ra
      -- 
    ra_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_0, ack => concat_CP_34_elements(475)); -- 
    -- CP-element group 476:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	474 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	545 
    -- CP-element group 476: marked-successors 
    -- CP-element group 476: 	182 
    -- CP-element group 476: 	222 
    -- CP-element group 476: 	243 
    -- CP-element group 476: 	264 
    -- CP-element group 476: 	474 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_update_completed_
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/$exit
      -- CP-element group 476: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1202_Update/ca
      -- 
    ca_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1202_inst_ack_1, ack => concat_CP_34_elements(476)); -- 
    -- CP-element group 477:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	386 
    -- CP-element group 477: 	394 
    -- CP-element group 477: 	398 
    -- CP-element group 477: marked-predecessors 
    -- CP-element group 477: 	479 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_sample_start_
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/$entry
      -- CP-element group 477: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/req
      -- 
    req_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(477), ack => W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_0); -- 
    concat_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(479);
      gj_concat_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: marked-predecessors 
    -- CP-element group 478: 	480 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	480 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_update_start_
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/req
      -- 
    req_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(478), ack => W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_1); -- 
    concat_cp_element_group_478: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_478"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(480);
      gj_concat_cp_element_group_478 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(478), clk => clk, reset => reset); --
    end block;
    -- CP-element group 479:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: successors 
    -- CP-element group 479: marked-successors 
    -- CP-element group 479: 	384 
    -- CP-element group 479: 	392 
    -- CP-element group 479: 	396 
    -- CP-element group 479: 	477 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_sample_completed_
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/$exit
      -- CP-element group 479: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Sample/ack
      -- 
    ack_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_0, ack => concat_CP_34_elements(479)); -- 
    -- CP-element group 480:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	551 
    -- CP-element group 480: marked-successors 
    -- CP-element group 480: 	478 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_update_completed_
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/$exit
      -- CP-element group 480: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1206_Update/ack
      -- 
    ack_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_1, ack => concat_CP_34_elements(480)); -- 
    -- CP-element group 481:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	386 
    -- CP-element group 481: 	394 
    -- CP-element group 481: 	398 
    -- CP-element group 481: marked-predecessors 
    -- CP-element group 481: 	483 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	483 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/req
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_sample_start_
      -- 
    req_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(481), ack => W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_0); -- 
    concat_cp_element_group_481: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_481"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(483);
      gj_concat_cp_element_group_481 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(481), clk => clk, reset => reset); --
    end block;
    -- CP-element group 482:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	179 
    -- CP-element group 482: marked-predecessors 
    -- CP-element group 482: 	484 
    -- CP-element group 482: 	547 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	484 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/req
      -- CP-element group 482: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_update_start_
      -- 
    req_2568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(482), ack => W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_1); -- 
    concat_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(484) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	481 
    -- CP-element group 483: successors 
    -- CP-element group 483: marked-successors 
    -- CP-element group 483: 	384 
    -- CP-element group 483: 	392 
    -- CP-element group 483: 	396 
    -- CP-element group 483: 	481 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/ack
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_sample_completed_
      -- 
    ack_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_0, ack => concat_CP_34_elements(483)); -- 
    -- CP-element group 484:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	545 
    -- CP-element group 484: marked-successors 
    -- CP-element group 484: 	182 
    -- CP-element group 484: 	222 
    -- CP-element group 484: 	243 
    -- CP-element group 484: 	264 
    -- CP-element group 484: 	482 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_Update/ack
      -- CP-element group 484: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1215_update_completed_
      -- 
    ack_2569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_1, ack => concat_CP_34_elements(484)); -- 
    -- CP-element group 485:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	386 
    -- CP-element group 485: 	394 
    -- CP-element group 485: 	398 
    -- CP-element group 485: marked-predecessors 
    -- CP-element group 485: 	487 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	487 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/req
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/$entry
      -- CP-element group 485: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_sample_start_
      -- 
    req_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(485), ack => W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_0); -- 
    concat_cp_element_group_485: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_485"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(487);
      gj_concat_cp_element_group_485 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(485), clk => clk, reset => reset); --
    end block;
    -- CP-element group 486:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	179 
    -- CP-element group 486: marked-predecessors 
    -- CP-element group 486: 	488 
    -- CP-element group 486: 	547 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	488 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/req
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/$entry
      -- CP-element group 486: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_update_start_
      -- 
    req_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(486), ack => W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_1); -- 
    concat_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(488) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	485 
    -- CP-element group 487: successors 
    -- CP-element group 487: marked-successors 
    -- CP-element group 487: 	384 
    -- CP-element group 487: 	392 
    -- CP-element group 487: 	396 
    -- CP-element group 487: 	485 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/ack
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_sample_completed_
      -- 
    ack_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_0, ack => concat_CP_34_elements(487)); -- 
    -- CP-element group 488:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	486 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	545 
    -- CP-element group 488: marked-successors 
    -- CP-element group 488: 	182 
    -- CP-element group 488: 	222 
    -- CP-element group 488: 	243 
    -- CP-element group 488: 	264 
    -- CP-element group 488: 	486 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/assign_stmt_1223_Update/ack
      -- 
    ack_2583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_1, ack => concat_CP_34_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	386 
    -- CP-element group 489: 	394 
    -- CP-element group 489: 	398 
    -- CP-element group 489: 	456 
    -- CP-element group 489: 	468 
    -- CP-element group 489: marked-predecessors 
    -- CP-element group 489: 	491 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	491 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/rr
      -- 
    rr_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(489), ack => type_cast_1238_inst_req_0); -- 
    concat_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(456) & concat_CP_34_elements(468) & concat_CP_34_elements(491);
      gj_concat_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	179 
    -- CP-element group 490: marked-predecessors 
    -- CP-element group 490: 	492 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	492 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/cr
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_update_start_
      -- CP-element group 490: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/$entry
      -- 
    cr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(490), ack => type_cast_1238_inst_req_1); -- 
    concat_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(492);
      gj_concat_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	489 
    -- CP-element group 491: successors 
    -- CP-element group 491: marked-successors 
    -- CP-element group 491: 	384 
    -- CP-element group 491: 	392 
    -- CP-element group 491: 	396 
    -- CP-element group 491: 	454 
    -- CP-element group 491: 	466 
    -- CP-element group 491: 	489 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Sample/ra
      -- 
    ra_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => concat_CP_34_elements(491)); -- 
    -- CP-element group 492:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	490 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	551 
    -- CP-element group 492: marked-successors 
    -- CP-element group 492: 	222 
    -- CP-element group 492: 	490 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/ca
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1238_update_completed_
      -- 
    ca_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => concat_CP_34_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	386 
    -- CP-element group 493: 	394 
    -- CP-element group 493: 	398 
    -- CP-element group 493: 	456 
    -- CP-element group 493: 	468 
    -- CP-element group 493: marked-predecessors 
    -- CP-element group 493: 	495 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	495 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_sample_start_
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/$entry
      -- CP-element group 493: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/rr
      -- 
    rr_2605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(493), ack => type_cast_1242_inst_req_0); -- 
    concat_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(456) & concat_CP_34_elements(468) & concat_CP_34_elements(495);
      gj_concat_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	179 
    -- CP-element group 494: marked-predecessors 
    -- CP-element group 494: 	496 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	496 
    -- CP-element group 494:  members (3) 
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_update_start_
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/$entry
      -- CP-element group 494: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/cr
      -- 
    cr_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(494), ack => type_cast_1242_inst_req_1); -- 
    concat_cp_element_group_494: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_494"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(496);
      gj_concat_cp_element_group_494 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(494), clk => clk, reset => reset); --
    end block;
    -- CP-element group 495:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	493 
    -- CP-element group 495: successors 
    -- CP-element group 495: marked-successors 
    -- CP-element group 495: 	384 
    -- CP-element group 495: 	392 
    -- CP-element group 495: 	396 
    -- CP-element group 495: 	454 
    -- CP-element group 495: 	466 
    -- CP-element group 495: 	493 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_sample_completed_
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/$exit
      -- CP-element group 495: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Sample/ra
      -- 
    ra_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_0, ack => concat_CP_34_elements(495)); -- 
    -- CP-element group 496:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	494 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	551 
    -- CP-element group 496: marked-successors 
    -- CP-element group 496: 	222 
    -- CP-element group 496: 	494 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/$exit
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_update_completed_
      -- CP-element group 496: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1242_Update/ca
      -- 
    ca_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1242_inst_ack_1, ack => concat_CP_34_elements(496)); -- 
    -- CP-element group 497:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	227 
    -- CP-element group 497: marked-predecessors 
    -- CP-element group 497: 	499 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	499 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_sample_start_
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/rr
      -- CP-element group 497: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/$entry
      -- 
    rr_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(497), ack => type_cast_1246_inst_req_0); -- 
    concat_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(227) & concat_CP_34_elements(499);
      gj_concat_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: marked-predecessors 
    -- CP-element group 498: 	500 
    -- CP-element group 498: 	503 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	500 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/cr
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/$entry
      -- CP-element group 498: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_update_start_
      -- 
    cr_2624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(498), ack => type_cast_1246_inst_req_1); -- 
    concat_cp_element_group_498: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_498"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(500) & concat_CP_34_elements(503);
      gj_concat_cp_element_group_498 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 499:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	497 
    -- CP-element group 499: successors 
    -- CP-element group 499: marked-successors 
    -- CP-element group 499: 	223 
    -- CP-element group 499: 	497 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/ra
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Sample/$exit
      -- CP-element group 499: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_sample_completed_
      -- 
    ra_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_0, ack => concat_CP_34_elements(499)); -- 
    -- CP-element group 500:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	498 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500: marked-successors 
    -- CP-element group 500: 	498 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/ca
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_Update/$exit
      -- CP-element group 500: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1246_update_completed_
      -- 
    ca_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_1, ack => concat_CP_34_elements(500)); -- 
    -- CP-element group 501:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	366 
    -- CP-element group 501: 	378 
    -- CP-element group 501: 	500 
    -- CP-element group 501: marked-predecessors 
    -- CP-element group 501: 	503 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	503 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/req
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/$entry
      -- CP-element group 501: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_sample_start_
      -- 
    req_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(501), ack => MUX_1253_inst_req_0); -- 
    concat_cp_element_group_501: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_501"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(378) & concat_CP_34_elements(500) & concat_CP_34_elements(503);
      gj_concat_cp_element_group_501 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(501), clk => clk, reset => reset); --
    end block;
    -- CP-element group 502:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	179 
    -- CP-element group 502: marked-predecessors 
    -- CP-element group 502: 	504 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	504 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/req
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_update_start_
      -- CP-element group 502: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/$entry
      -- 
    req_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(502), ack => MUX_1253_inst_req_1); -- 
    concat_cp_element_group_502: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_502"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(504);
      gj_concat_cp_element_group_502 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(502), clk => clk, reset => reset); --
    end block;
    -- CP-element group 503:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	501 
    -- CP-element group 503: successors 
    -- CP-element group 503: marked-successors 
    -- CP-element group 503: 	364 
    -- CP-element group 503: 	376 
    -- CP-element group 503: 	498 
    -- CP-element group 503: 	501 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/ack
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_start/$exit
      -- CP-element group 503: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_sample_completed_
      -- 
    ack_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1253_inst_ack_0, ack => concat_CP_34_elements(503)); -- 
    -- CP-element group 504:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	502 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	551 
    -- CP-element group 504: marked-successors 
    -- CP-element group 504: 	222 
    -- CP-element group 504: 	502 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/$exit
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_update_completed_
      -- CP-element group 504: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1253_complete/ack
      -- 
    ack_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1253_inst_ack_1, ack => concat_CP_34_elements(504)); -- 
    -- CP-element group 505:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	386 
    -- CP-element group 505: 	394 
    -- CP-element group 505: 	398 
    -- CP-element group 505: 	460 
    -- CP-element group 505: 	464 
    -- CP-element group 505: marked-predecessors 
    -- CP-element group 505: 	507 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	507 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_sample_start_
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/$entry
      -- CP-element group 505: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/rr
      -- 
    rr_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(505), ack => type_cast_1266_inst_req_0); -- 
    concat_cp_element_group_505: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_505"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(460) & concat_CP_34_elements(464) & concat_CP_34_elements(507);
      gj_concat_cp_element_group_505 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(505), clk => clk, reset => reset); --
    end block;
    -- CP-element group 506:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	179 
    -- CP-element group 506: marked-predecessors 
    -- CP-element group 506: 	508 
    -- CP-element group 506: 	547 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	508 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_update_start_
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/$entry
      -- CP-element group 506: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/cr
      -- 
    cr_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(506), ack => type_cast_1266_inst_req_1); -- 
    concat_cp_element_group_506: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_506"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(508) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_506 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(506), clk => clk, reset => reset); --
    end block;
    -- CP-element group 507:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	505 
    -- CP-element group 507: successors 
    -- CP-element group 507: marked-successors 
    -- CP-element group 507: 	384 
    -- CP-element group 507: 	392 
    -- CP-element group 507: 	396 
    -- CP-element group 507: 	458 
    -- CP-element group 507: 	462 
    -- CP-element group 507: 	505 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_sample_completed_
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/$exit
      -- CP-element group 507: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Sample/ra
      -- 
    ra_2648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => concat_CP_34_elements(507)); -- 
    -- CP-element group 508:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	506 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	545 
    -- CP-element group 508: marked-successors 
    -- CP-element group 508: 	182 
    -- CP-element group 508: 	506 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_update_completed_
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/$exit
      -- CP-element group 508: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1266_Update/ca
      -- 
    ca_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => concat_CP_34_elements(508)); -- 
    -- CP-element group 509:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	386 
    -- CP-element group 509: 	394 
    -- CP-element group 509: 	398 
    -- CP-element group 509: 	460 
    -- CP-element group 509: 	464 
    -- CP-element group 509: marked-predecessors 
    -- CP-element group 509: 	511 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	511 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/rr
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/$entry
      -- CP-element group 509: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_sample_start_
      -- 
    rr_2661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(509), ack => type_cast_1270_inst_req_0); -- 
    concat_cp_element_group_509: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_509"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(460) & concat_CP_34_elements(464) & concat_CP_34_elements(511);
      gj_concat_cp_element_group_509 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(509), clk => clk, reset => reset); --
    end block;
    -- CP-element group 510:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	179 
    -- CP-element group 510: marked-predecessors 
    -- CP-element group 510: 	512 
    -- CP-element group 510: 	547 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/$entry
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/cr
      -- CP-element group 510: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_update_start_
      -- 
    cr_2666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(510), ack => type_cast_1270_inst_req_1); -- 
    concat_cp_element_group_510: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_510"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(512) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_510 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(510), clk => clk, reset => reset); --
    end block;
    -- CP-element group 511:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	509 
    -- CP-element group 511: successors 
    -- CP-element group 511: marked-successors 
    -- CP-element group 511: 	384 
    -- CP-element group 511: 	392 
    -- CP-element group 511: 	396 
    -- CP-element group 511: 	458 
    -- CP-element group 511: 	462 
    -- CP-element group 511: 	509 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/ra
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Sample/$exit
      -- CP-element group 511: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_sample_completed_
      -- 
    ra_2662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_0, ack => concat_CP_34_elements(511)); -- 
    -- CP-element group 512:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	545 
    -- CP-element group 512: marked-successors 
    -- CP-element group 512: 	182 
    -- CP-element group 512: 	510 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/ca
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_Update/$exit
      -- CP-element group 512: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1270_update_completed_
      -- 
    ca_2667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_1, ack => concat_CP_34_elements(512)); -- 
    -- CP-element group 513:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	288 
    -- CP-element group 513: 	350 
    -- CP-element group 513: 	354 
    -- CP-element group 513: marked-predecessors 
    -- CP-element group 513: 	515 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	515 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_sample_start_
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/rr
      -- CP-element group 513: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/$entry
      -- 
    rr_2675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(513), ack => type_cast_1274_inst_req_0); -- 
    concat_cp_element_group_513: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_513"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(350) & concat_CP_34_elements(354) & concat_CP_34_elements(515);
      gj_concat_cp_element_group_513 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(513), clk => clk, reset => reset); --
    end block;
    -- CP-element group 514:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: marked-predecessors 
    -- CP-element group 514: 	516 
    -- CP-element group 514: 	519 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	516 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_update_start_
      -- 
    cr_2680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(514), ack => type_cast_1274_inst_req_1); -- 
    concat_cp_element_group_514: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_514"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(516) & concat_CP_34_elements(519);
      gj_concat_cp_element_group_514 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(514), clk => clk, reset => reset); --
    end block;
    -- CP-element group 515:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	513 
    -- CP-element group 515: successors 
    -- CP-element group 515: marked-successors 
    -- CP-element group 515: 	286 
    -- CP-element group 515: 	348 
    -- CP-element group 515: 	352 
    -- CP-element group 515: 	513 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/ra
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Sample/$exit
      -- CP-element group 515: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_sample_completed_
      -- 
    ra_2676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_0, ack => concat_CP_34_elements(515)); -- 
    -- CP-element group 516:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	514 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	517 
    -- CP-element group 516: marked-successors 
    -- CP-element group 516: 	514 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/ca
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_Update/$exit
      -- CP-element group 516: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1274_update_completed_
      -- 
    ca_2681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_1, ack => concat_CP_34_elements(516)); -- 
    -- CP-element group 517:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	366 
    -- CP-element group 517: 	378 
    -- CP-element group 517: 	516 
    -- CP-element group 517: marked-predecessors 
    -- CP-element group 517: 	519 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	519 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/req
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/$entry
      -- CP-element group 517: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_sample_start_
      -- 
    req_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(517), ack => MUX_1281_inst_req_0); -- 
    concat_cp_element_group_517: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_517"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(378) & concat_CP_34_elements(516) & concat_CP_34_elements(519);
      gj_concat_cp_element_group_517 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(517), clk => clk, reset => reset); --
    end block;
    -- CP-element group 518:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	179 
    -- CP-element group 518: marked-predecessors 
    -- CP-element group 518: 	520 
    -- CP-element group 518: 	547 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	520 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/req
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/$entry
      -- CP-element group 518: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_update_start_
      -- 
    req_2694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(518), ack => MUX_1281_inst_req_1); -- 
    concat_cp_element_group_518: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_518"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(520) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_518 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(518), clk => clk, reset => reset); --
    end block;
    -- CP-element group 519:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	517 
    -- CP-element group 519: successors 
    -- CP-element group 519: marked-successors 
    -- CP-element group 519: 	364 
    -- CP-element group 519: 	376 
    -- CP-element group 519: 	514 
    -- CP-element group 519: 	517 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/ack
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_start/$exit
      -- CP-element group 519: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_sample_completed_
      -- 
    ack_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1281_inst_ack_0, ack => concat_CP_34_elements(519)); -- 
    -- CP-element group 520:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	518 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	545 
    -- CP-element group 520: marked-successors 
    -- CP-element group 520: 	182 
    -- CP-element group 520: 	518 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/ack
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_complete/$exit
      -- CP-element group 520: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1281_update_completed_
      -- 
    ack_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1281_inst_ack_1, ack => concat_CP_34_elements(520)); -- 
    -- CP-element group 521:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	288 
    -- CP-element group 521: 	342 
    -- CP-element group 521: 	362 
    -- CP-element group 521: marked-predecessors 
    -- CP-element group 521: 	523 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	523 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/rr
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_sample_start_
      -- 
    rr_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(521), ack => type_cast_1294_inst_req_0); -- 
    concat_cp_element_group_521: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_521"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(342) & concat_CP_34_elements(362) & concat_CP_34_elements(523);
      gj_concat_cp_element_group_521 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(521), clk => clk, reset => reset); --
    end block;
    -- CP-element group 522:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	179 
    -- CP-element group 522: marked-predecessors 
    -- CP-element group 522: 	524 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	524 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/cr
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/$entry
      -- CP-element group 522: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_update_start_
      -- 
    cr_2708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(522), ack => type_cast_1294_inst_req_1); -- 
    concat_cp_element_group_522: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_522"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(524);
      gj_concat_cp_element_group_522 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(522), clk => clk, reset => reset); --
    end block;
    -- CP-element group 523:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	521 
    -- CP-element group 523: successors 
    -- CP-element group 523: marked-successors 
    -- CP-element group 523: 	286 
    -- CP-element group 523: 	340 
    -- CP-element group 523: 	360 
    -- CP-element group 523: 	521 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/ra
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_sample_completed_
      -- 
    ra_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_0, ack => concat_CP_34_elements(523)); -- 
    -- CP-element group 524:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	522 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	551 
    -- CP-element group 524: marked-successors 
    -- CP-element group 524: 	243 
    -- CP-element group 524: 	522 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/ca
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1294_update_completed_
      -- 
    ca_2709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1294_inst_ack_1, ack => concat_CP_34_elements(524)); -- 
    -- CP-element group 525:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	288 
    -- CP-element group 525: 	342 
    -- CP-element group 525: 	362 
    -- CP-element group 525: marked-predecessors 
    -- CP-element group 525: 	527 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	527 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/rr
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/$entry
      -- CP-element group 525: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_sample_start_
      -- 
    rr_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(525), ack => type_cast_1298_inst_req_0); -- 
    concat_cp_element_group_525: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_525"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(288) & concat_CP_34_elements(342) & concat_CP_34_elements(362) & concat_CP_34_elements(527);
      gj_concat_cp_element_group_525 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(525), clk => clk, reset => reset); --
    end block;
    -- CP-element group 526:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: marked-predecessors 
    -- CP-element group 526: 	528 
    -- CP-element group 526: 	531 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	528 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/cr
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/$entry
      -- CP-element group 526: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_update_start_
      -- 
    cr_2722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(526), ack => type_cast_1298_inst_req_1); -- 
    concat_cp_element_group_526: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_526"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(528) & concat_CP_34_elements(531);
      gj_concat_cp_element_group_526 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(526), clk => clk, reset => reset); --
    end block;
    -- CP-element group 527:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	525 
    -- CP-element group 527: successors 
    -- CP-element group 527: marked-successors 
    -- CP-element group 527: 	286 
    -- CP-element group 527: 	340 
    -- CP-element group 527: 	360 
    -- CP-element group 527: 	525 
    -- CP-element group 527:  members (3) 
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/ra
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Sample/$exit
      -- CP-element group 527: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_sample_completed_
      -- 
    ra_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_0, ack => concat_CP_34_elements(527)); -- 
    -- CP-element group 528:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	526 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528: marked-successors 
    -- CP-element group 528: 	526 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/ca
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_Update/$exit
      -- CP-element group 528: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1298_update_completed_
      -- 
    ca_2723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_1, ack => concat_CP_34_elements(528)); -- 
    -- CP-element group 529:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	366 
    -- CP-element group 529: 	378 
    -- CP-element group 529: 	528 
    -- CP-element group 529: marked-predecessors 
    -- CP-element group 529: 	531 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	531 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_sample_start_
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/req
      -- CP-element group 529: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/$entry
      -- 
    req_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(529), ack => MUX_1305_inst_req_0); -- 
    concat_cp_element_group_529: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_529"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(378) & concat_CP_34_elements(528) & concat_CP_34_elements(531);
      gj_concat_cp_element_group_529 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(529), clk => clk, reset => reset); --
    end block;
    -- CP-element group 530:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	179 
    -- CP-element group 530: marked-predecessors 
    -- CP-element group 530: 	532 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/$entry
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/req
      -- CP-element group 530: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_update_start_
      -- 
    req_2736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(530), ack => MUX_1305_inst_req_1); -- 
    concat_cp_element_group_530: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_530"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(532);
      gj_concat_cp_element_group_530 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(530), clk => clk, reset => reset); --
    end block;
    -- CP-element group 531:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	529 
    -- CP-element group 531: successors 
    -- CP-element group 531: marked-successors 
    -- CP-element group 531: 	364 
    -- CP-element group 531: 	376 
    -- CP-element group 531: 	526 
    -- CP-element group 531: 	529 
    -- CP-element group 531:  members (3) 
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/ack
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_sample_completed_
      -- CP-element group 531: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_start/$exit
      -- 
    ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1305_inst_ack_0, ack => concat_CP_34_elements(531)); -- 
    -- CP-element group 532:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	551 
    -- CP-element group 532: marked-successors 
    -- CP-element group 532: 	243 
    -- CP-element group 532: 	530 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/$exit
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_complete/ack
      -- CP-element group 532: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1305_update_completed_
      -- 
    ack_2737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1305_inst_ack_1, ack => concat_CP_34_elements(532)); -- 
    -- CP-element group 533:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	386 
    -- CP-element group 533: 	394 
    -- CP-element group 533: 	398 
    -- CP-element group 533: 	452 
    -- CP-element group 533: 	472 
    -- CP-element group 533: marked-predecessors 
    -- CP-element group 533: 	535 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	535 
    -- CP-element group 533:  members (3) 
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_sample_start_
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/rr
      -- CP-element group 533: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/$entry
      -- 
    rr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(533), ack => type_cast_1320_inst_req_0); -- 
    concat_cp_element_group_533: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_533"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= concat_CP_34_elements(386) & concat_CP_34_elements(394) & concat_CP_34_elements(398) & concat_CP_34_elements(452) & concat_CP_34_elements(472) & concat_CP_34_elements(535);
      gj_concat_cp_element_group_533 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(533), clk => clk, reset => reset); --
    end block;
    -- CP-element group 534:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	179 
    -- CP-element group 534: marked-predecessors 
    -- CP-element group 534: 	536 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	536 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_update_start_
      -- 
    cr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(534), ack => type_cast_1320_inst_req_1); -- 
    concat_cp_element_group_534: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_534"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(536);
      gj_concat_cp_element_group_534 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(534), clk => clk, reset => reset); --
    end block;
    -- CP-element group 535:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	533 
    -- CP-element group 535: successors 
    -- CP-element group 535: marked-successors 
    -- CP-element group 535: 	384 
    -- CP-element group 535: 	392 
    -- CP-element group 535: 	396 
    -- CP-element group 535: 	450 
    -- CP-element group 535: 	470 
    -- CP-element group 535: 	533 
    -- CP-element group 535:  members (3) 
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_sample_completed_
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/ra
      -- CP-element group 535: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Sample/$exit
      -- 
    ra_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => concat_CP_34_elements(535)); -- 
    -- CP-element group 536:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	534 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	551 
    -- CP-element group 536: marked-successors 
    -- CP-element group 536: 	264 
    -- CP-element group 536: 	534 
    -- CP-element group 536:  members (3) 
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/ca
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_Update/$exit
      -- CP-element group 536: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1320_update_completed_
      -- 
    ca_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => concat_CP_34_elements(536)); -- 
    -- CP-element group 537:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	269 
    -- CP-element group 537: marked-predecessors 
    -- CP-element group 537: 	539 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	539 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_sample_start_
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/$entry
      -- CP-element group 537: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/rr
      -- 
    rr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(537), ack => type_cast_1324_inst_req_0); -- 
    concat_cp_element_group_537: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_537"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(269) & concat_CP_34_elements(539);
      gj_concat_cp_element_group_537 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(537), clk => clk, reset => reset); --
    end block;
    -- CP-element group 538:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: marked-predecessors 
    -- CP-element group 538: 	540 
    -- CP-element group 538: 	543 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	540 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/cr
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_update_start_
      -- CP-element group 538: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/$entry
      -- 
    cr_2764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(538), ack => type_cast_1324_inst_req_1); -- 
    concat_cp_element_group_538: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_538"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(540) & concat_CP_34_elements(543);
      gj_concat_cp_element_group_538 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(538), clk => clk, reset => reset); --
    end block;
    -- CP-element group 539:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	537 
    -- CP-element group 539: successors 
    -- CP-element group 539: marked-successors 
    -- CP-element group 539: 	265 
    -- CP-element group 539: 	537 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Sample/ra
      -- 
    ra_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1324_inst_ack_0, ack => concat_CP_34_elements(539)); -- 
    -- CP-element group 540:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	538 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540: marked-successors 
    -- CP-element group 540: 	538 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1324_Update/ca
      -- 
    ca_2765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1324_inst_ack_1, ack => concat_CP_34_elements(540)); -- 
    -- CP-element group 541:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	366 
    -- CP-element group 541: 	378 
    -- CP-element group 541: 	540 
    -- CP-element group 541: marked-predecessors 
    -- CP-element group 541: 	543 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	543 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/req
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_sample_start_
      -- CP-element group 541: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/$entry
      -- 
    req_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(541), ack => MUX_1331_inst_req_0); -- 
    concat_cp_element_group_541: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_541"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_CP_34_elements(366) & concat_CP_34_elements(378) & concat_CP_34_elements(540) & concat_CP_34_elements(543);
      gj_concat_cp_element_group_541 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(541), clk => clk, reset => reset); --
    end block;
    -- CP-element group 542:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	179 
    -- CP-element group 542: marked-predecessors 
    -- CP-element group 542: 	544 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	544 
    -- CP-element group 542:  members (3) 
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/req
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/$entry
      -- CP-element group 542: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_update_start_
      -- 
    req_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(542), ack => MUX_1331_inst_req_1); -- 
    concat_cp_element_group_542: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_542"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(179) & concat_CP_34_elements(544);
      gj_concat_cp_element_group_542 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(542), clk => clk, reset => reset); --
    end block;
    -- CP-element group 543:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	541 
    -- CP-element group 543: successors 
    -- CP-element group 543: marked-successors 
    -- CP-element group 543: 	364 
    -- CP-element group 543: 	376 
    -- CP-element group 543: 	538 
    -- CP-element group 543: 	541 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/ack
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_start/$exit
      -- CP-element group 543: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_sample_completed_
      -- 
    ack_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1331_inst_ack_0, ack => concat_CP_34_elements(543)); -- 
    -- CP-element group 544:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	542 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	551 
    -- CP-element group 544: marked-successors 
    -- CP-element group 544: 	264 
    -- CP-element group 544: 	542 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/ack
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_complete/$exit
      -- CP-element group 544: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/MUX_1331_update_completed_
      -- 
    ack_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1331_inst_ack_1, ack => concat_CP_34_elements(544)); -- 
    -- CP-element group 545:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	476 
    -- CP-element group 545: 	484 
    -- CP-element group 545: 	488 
    -- CP-element group 545: 	508 
    -- CP-element group 545: 	512 
    -- CP-element group 545: 	520 
    -- CP-element group 545: marked-predecessors 
    -- CP-element group 545: 	547 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	547 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_sample_start_
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/rr
      -- CP-element group 545: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/$entry
      -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(545), ack => type_cast_1346_inst_req_0); -- 
    concat_cp_element_group_545: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 27) := "concat_cp_element_group_545"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= concat_CP_34_elements(476) & concat_CP_34_elements(484) & concat_CP_34_elements(488) & concat_CP_34_elements(508) & concat_CP_34_elements(512) & concat_CP_34_elements(520) & concat_CP_34_elements(547);
      gj_concat_cp_element_group_545 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(545), clk => clk, reset => reset); --
    end block;
    -- CP-element group 546:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: marked-predecessors 
    -- CP-element group 546: 	548 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	548 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/cr
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/$entry
      -- CP-element group 546: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_update_start_
      -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(546), ack => type_cast_1346_inst_req_1); -- 
    concat_cp_element_group_546: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_546"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_CP_34_elements(548);
      gj_concat_cp_element_group_546 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(546), clk => clk, reset => reset); --
    end block;
    -- CP-element group 547:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	545 
    -- CP-element group 547: successors 
    -- CP-element group 547: marked-successors 
    -- CP-element group 547: 	474 
    -- CP-element group 547: 	482 
    -- CP-element group 547: 	486 
    -- CP-element group 547: 	506 
    -- CP-element group 547: 	510 
    -- CP-element group 547: 	518 
    -- CP-element group 547: 	545 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/ra
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_sample_completed_
      -- CP-element group 547: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Sample/$exit
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => concat_CP_34_elements(547)); -- 
    -- CP-element group 548:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	546 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	177 
    -- CP-element group 548: marked-successors 
    -- CP-element group 548: 	546 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/ca
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_Update/$exit
      -- CP-element group 548: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/type_cast_1346_update_completed_
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => concat_CP_34_elements(548)); -- 
    -- CP-element group 549:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	176 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	177 
    -- CP-element group 549:  members (1) 
      -- CP-element group 549: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_CP_34_elements(549) is a control-delay.
    cp_element_549_delay: control_delay_element  generic map(name => " 549_delay", delay_value => 1)  port map(req => concat_CP_34_elements(176), ack => concat_CP_34_elements(549), clk => clk, reset =>reset);
    -- CP-element group 550:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	337 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	445 
    -- CP-element group 550:  members (1) 
      -- CP-element group 550: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/ptr_deref_910_ptr_deref_1113_delay
      -- 
    -- Element group concat_CP_34_elements(550) is a control-delay.
    cp_element_550_delay: control_delay_element  generic map(name => " 550_delay", delay_value => 1)  port map(req => concat_CP_34_elements(337), ack => concat_CP_34_elements(550), clk => clk, reset =>reset);
    -- CP-element group 551:  join  transition  bypass  pipeline-parent 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	300 
    -- CP-element group 551: 	323 
    -- CP-element group 551: 	330 
    -- CP-element group 551: 	338 
    -- CP-element group 551: 	346 
    -- CP-element group 551: 	358 
    -- CP-element group 551: 	370 
    -- CP-element group 551: 	390 
    -- CP-element group 551: 	410 
    -- CP-element group 551: 	433 
    -- CP-element group 551: 	440 
    -- CP-element group 551: 	447 
    -- CP-element group 551: 	448 
    -- CP-element group 551: 	480 
    -- CP-element group 551: 	492 
    -- CP-element group 551: 	496 
    -- CP-element group 551: 	504 
    -- CP-element group 551: 	524 
    -- CP-element group 551: 	532 
    -- CP-element group 551: 	536 
    -- CP-element group 551: 	544 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	173 
    -- CP-element group 551:  members (1) 
      -- CP-element group 551: 	 branch_block_stmt_23/do_while_stmt_817/do_while_stmt_817_loop_body/$exit
      -- 
    concat_cp_element_group_551: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_551"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= concat_CP_34_elements(300) & concat_CP_34_elements(323) & concat_CP_34_elements(330) & concat_CP_34_elements(338) & concat_CP_34_elements(346) & concat_CP_34_elements(358) & concat_CP_34_elements(370) & concat_CP_34_elements(390) & concat_CP_34_elements(410) & concat_CP_34_elements(433) & concat_CP_34_elements(440) & concat_CP_34_elements(447) & concat_CP_34_elements(448) & concat_CP_34_elements(480) & concat_CP_34_elements(492) & concat_CP_34_elements(496) & concat_CP_34_elements(504) & concat_CP_34_elements(524) & concat_CP_34_elements(532) & concat_CP_34_elements(536) & concat_CP_34_elements(544);
      gj_concat_cp_element_group_551 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 552:  transition  input  bypass  pipeline-parent 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	172 
    -- CP-element group 552: successors 
    -- CP-element group 552:  members (2) 
      -- CP-element group 552: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/ack
      -- CP-element group 552: 	 branch_block_stmt_23/do_while_stmt_817/loop_exit/$exit
      -- 
    ack_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_817_branch_ack_0, ack => concat_CP_34_elements(552)); -- 
    -- CP-element group 553:  transition  input  bypass  pipeline-parent 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	172 
    -- CP-element group 553: successors 
    -- CP-element group 553:  members (2) 
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/$exit
      -- CP-element group 553: 	 branch_block_stmt_23/do_while_stmt_817/loop_taken/ack
      -- 
    ack_2804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_817_branch_ack_1, ack => concat_CP_34_elements(553)); -- 
    -- CP-element group 554:  transition  bypass  pipeline-parent 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	170 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	1 
    -- CP-element group 554:  members (1) 
      -- CP-element group 554: 	 branch_block_stmt_23/do_while_stmt_817/$exit
      -- 
    concat_CP_34_elements(554) <= concat_CP_34_elements(170);
    -- CP-element group 555:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	1 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	557 
    -- CP-element group 555: 	558 
    -- CP-element group 555:  members (18) 
      -- CP-element group 555: 	 branch_block_stmt_23/merge_stmt_1363__exit__
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369__entry__
      -- CP-element group 555: 	 branch_block_stmt_23/ifx_xend300_whilex_xend_PhiReq/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/merge_stmt_1363_PhiReqMerge
      -- CP-element group 555: 	 branch_block_stmt_23/ifx_xend300_whilex_xend_PhiReq/$exit
      -- CP-element group 555: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/$exit
      -- CP-element group 555: 	 branch_block_stmt_23/merge_stmt_1363_PhiAck/dummy
      -- CP-element group 555: 	 branch_block_stmt_23/if_stmt_1359_if_link/$exit
      -- CP-element group 555: 	 branch_block_stmt_23/if_stmt_1359_if_link/if_choice_transition
      -- CP-element group 555: 	 branch_block_stmt_23/ifx_xend300_whilex_xend
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_sample_start_
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_update_start_
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/rr
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/$entry
      -- CP-element group 555: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/cr
      -- 
    if_choice_transition_2818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 555_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_1, ack => concat_CP_34_elements(555)); -- 
    rr_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(555), ack => type_cast_1368_inst_req_0); -- 
    cr_2839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(555), ack => type_cast_1368_inst_req_1); -- 
    -- CP-element group 556:  merge  transition  place  input  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	1 
    -- CP-element group 556: successors 
    -- CP-element group 556:  members (5) 
      -- CP-element group 556: 	 branch_block_stmt_23/if_stmt_1359__exit__
      -- CP-element group 556: 	 branch_block_stmt_23/merge_stmt_1363__entry__
      -- CP-element group 556: 	 branch_block_stmt_23/merge_stmt_1363_dead_link/$entry
      -- CP-element group 556: 	 branch_block_stmt_23/if_stmt_1359_else_link/$exit
      -- CP-element group 556: 	 branch_block_stmt_23/if_stmt_1359_else_link/else_choice_transition
      -- 
    else_choice_transition_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1359_branch_ack_0, ack => concat_CP_34_elements(556)); -- 
    -- CP-element group 557:  transition  input  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	555 
    -- CP-element group 557: successors 
    -- CP-element group 557:  members (3) 
      -- CP-element group 557: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_sample_completed_
      -- CP-element group 557: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/$exit
      -- CP-element group 557: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Sample/ra
      -- 
    ra_2835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => concat_CP_34_elements(557)); -- 
    -- CP-element group 558:  fork  transition  place  input  output  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	555 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	559 
    -- CP-element group 558: 	560 
    -- CP-element group 558: 	562 
    -- CP-element group 558: 	564 
    -- CP-element group 558: 	566 
    -- CP-element group 558: 	568 
    -- CP-element group 558: 	570 
    -- CP-element group 558: 	572 
    -- CP-element group 558: 	574 
    -- CP-element group 558: 	576 
    -- CP-element group 558: 	578 
    -- CP-element group 558:  members (40) 
      -- CP-element group 558: 	 branch_block_stmt_23/assign_stmt_1369__exit__
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480__entry__
      -- CP-element group 558: 	 branch_block_stmt_23/assign_stmt_1369/$exit
      -- CP-element group 558: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_update_completed_
      -- CP-element group 558: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/$exit
      -- CP-element group 558: 	 branch_block_stmt_23/assign_stmt_1369/type_cast_1368_Update/ca
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_sample_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/crr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/ccr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/cr
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_update_start_
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/$entry
      -- CP-element group 558: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/cr
      -- 
    ca_2840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 558_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => concat_CP_34_elements(558)); -- 
    crr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => call_stmt_1372_call_req_0); -- 
    ccr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => call_stmt_1372_call_req_1); -- 
    cr_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1376_inst_req_1); -- 
    cr_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1385_inst_req_1); -- 
    cr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1395_inst_req_1); -- 
    cr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1405_inst_req_1); -- 
    cr_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1415_inst_req_1); -- 
    cr_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1425_inst_req_1); -- 
    cr_2954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1435_inst_req_1); -- 
    cr_2968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1445_inst_req_1); -- 
    cr_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(558), ack => type_cast_1455_inst_req_1); -- 
    -- CP-element group 559:  transition  input  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	558 
    -- CP-element group 559: successors 
    -- CP-element group 559:  members (3) 
      -- CP-element group 559: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_sample_completed_
      -- CP-element group 559: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/$exit
      -- CP-element group 559: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Sample/cra
      -- 
    cra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1372_call_ack_0, ack => concat_CP_34_elements(559)); -- 
    -- CP-element group 560:  transition  input  output  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	558 
    -- CP-element group 560: successors 
    -- CP-element group 560: 	561 
    -- CP-element group 560:  members (6) 
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_update_completed_
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/$exit
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/call_stmt_1372_Update/cca
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_sample_start_
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/$entry
      -- CP-element group 560: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/rr
      -- 
    cca_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1372_call_ack_1, ack => concat_CP_34_elements(560)); -- 
    rr_2865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(560), ack => type_cast_1376_inst_req_0); -- 
    -- CP-element group 561:  transition  input  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	560 
    -- CP-element group 561: successors 
    -- CP-element group 561:  members (3) 
      -- CP-element group 561: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_sample_completed_
      -- CP-element group 561: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/$exit
      -- CP-element group 561: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Sample/ra
      -- 
    ra_2866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => concat_CP_34_elements(561)); -- 
    -- CP-element group 562:  fork  transition  input  output  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	558 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	563 
    -- CP-element group 562: 	565 
    -- CP-element group 562: 	567 
    -- CP-element group 562: 	569 
    -- CP-element group 562: 	571 
    -- CP-element group 562: 	573 
    -- CP-element group 562: 	575 
    -- CP-element group 562: 	577 
    -- CP-element group 562:  members (27) 
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_update_completed_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/$exit
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1376_Update/ca
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/rr
      -- 
    ca_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 562_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => concat_CP_34_elements(562)); -- 
    rr_2879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1385_inst_req_0); -- 
    rr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1395_inst_req_0); -- 
    rr_2907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1405_inst_req_0); -- 
    rr_2921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1415_inst_req_0); -- 
    rr_2935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1425_inst_req_0); -- 
    rr_2949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1435_inst_req_0); -- 
    rr_2963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1445_inst_req_0); -- 
    rr_2977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(562), ack => type_cast_1455_inst_req_0); -- 
    -- CP-element group 563:  transition  input  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	562 
    -- CP-element group 563: successors 
    -- CP-element group 563:  members (3) 
      -- CP-element group 563: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_sample_completed_
      -- CP-element group 563: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/$exit
      -- CP-element group 563: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Sample/ra
      -- 
    ra_2880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 563_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_0, ack => concat_CP_34_elements(563)); -- 
    -- CP-element group 564:  transition  input  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	558 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	599 
    -- CP-element group 564:  members (3) 
      -- CP-element group 564: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_update_completed_
      -- CP-element group 564: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/$exit
      -- CP-element group 564: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1385_Update/ca
      -- 
    ca_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_1, ack => concat_CP_34_elements(564)); -- 
    -- CP-element group 565:  transition  input  bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	562 
    -- CP-element group 565: successors 
    -- CP-element group 565:  members (3) 
      -- CP-element group 565: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_sample_completed_
      -- CP-element group 565: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/$exit
      -- CP-element group 565: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Sample/ra
      -- 
    ra_2894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => concat_CP_34_elements(565)); -- 
    -- CP-element group 566:  transition  input  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	558 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	596 
    -- CP-element group 566:  members (3) 
      -- CP-element group 566: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_update_completed_
      -- CP-element group 566: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/$exit
      -- CP-element group 566: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1395_Update/ca
      -- 
    ca_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_1, ack => concat_CP_34_elements(566)); -- 
    -- CP-element group 567:  transition  input  bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	562 
    -- CP-element group 567: successors 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_sample_completed_
      -- CP-element group 567: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/$exit
      -- CP-element group 567: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Sample/ra
      -- 
    ra_2908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_0, ack => concat_CP_34_elements(567)); -- 
    -- CP-element group 568:  transition  input  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	558 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	593 
    -- CP-element group 568:  members (3) 
      -- CP-element group 568: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_update_completed_
      -- CP-element group 568: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/$exit
      -- CP-element group 568: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1405_Update/ca
      -- 
    ca_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_1, ack => concat_CP_34_elements(568)); -- 
    -- CP-element group 569:  transition  input  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	562 
    -- CP-element group 569: successors 
    -- CP-element group 569:  members (3) 
      -- CP-element group 569: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_sample_completed_
      -- CP-element group 569: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/$exit
      -- CP-element group 569: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Sample/ra
      -- 
    ra_2922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_0, ack => concat_CP_34_elements(569)); -- 
    -- CP-element group 570:  transition  input  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	558 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	590 
    -- CP-element group 570:  members (3) 
      -- CP-element group 570: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_update_completed_
      -- CP-element group 570: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/$exit
      -- CP-element group 570: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1415_Update/ca
      -- 
    ca_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 570_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1415_inst_ack_1, ack => concat_CP_34_elements(570)); -- 
    -- CP-element group 571:  transition  input  bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	562 
    -- CP-element group 571: successors 
    -- CP-element group 571:  members (3) 
      -- CP-element group 571: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/$exit
      -- CP-element group 571: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Sample/ra
      -- 
    ra_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => concat_CP_34_elements(571)); -- 
    -- CP-element group 572:  transition  input  bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	558 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	587 
    -- CP-element group 572:  members (3) 
      -- CP-element group 572: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/$exit
      -- CP-element group 572: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1425_Update/ca
      -- 
    ca_2941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => concat_CP_34_elements(572)); -- 
    -- CP-element group 573:  transition  input  bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	562 
    -- CP-element group 573: successors 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_sample_completed_
      -- CP-element group 573: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/$exit
      -- CP-element group 573: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Sample/ra
      -- 
    ra_2950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_0, ack => concat_CP_34_elements(573)); -- 
    -- CP-element group 574:  transition  input  bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	558 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	584 
    -- CP-element group 574:  members (3) 
      -- CP-element group 574: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_update_completed_
      -- CP-element group 574: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/$exit
      -- CP-element group 574: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1435_Update/ca
      -- 
    ca_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1435_inst_ack_1, ack => concat_CP_34_elements(574)); -- 
    -- CP-element group 575:  transition  input  bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	562 
    -- CP-element group 575: successors 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_sample_completed_
      -- CP-element group 575: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/$exit
      -- CP-element group 575: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Sample/ra
      -- 
    ra_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_0, ack => concat_CP_34_elements(575)); -- 
    -- CP-element group 576:  transition  input  bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	558 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	581 
    -- CP-element group 576:  members (3) 
      -- CP-element group 576: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_update_completed_
      -- CP-element group 576: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/$exit
      -- CP-element group 576: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1445_Update/ca
      -- 
    ca_2969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1445_inst_ack_1, ack => concat_CP_34_elements(576)); -- 
    -- CP-element group 577:  transition  input  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	562 
    -- CP-element group 577: successors 
    -- CP-element group 577:  members (3) 
      -- CP-element group 577: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_sample_completed_
      -- CP-element group 577: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/$exit
      -- CP-element group 577: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Sample/ra
      -- 
    ra_2978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 577_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_0, ack => concat_CP_34_elements(577)); -- 
    -- CP-element group 578:  transition  input  output  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	558 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	579 
    -- CP-element group 578:  members (6) 
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_update_completed_
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/$exit
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/type_cast_1455_Update/ca
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_sample_start_
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/$entry
      -- CP-element group 578: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/req
      -- 
    ca_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 578_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1455_inst_ack_1, ack => concat_CP_34_elements(578)); -- 
    req_2991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(578), ack => WPIPE_Concat_output_pipe_1457_inst_req_0); -- 
    -- CP-element group 579:  transition  input  output  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	578 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	580 
    -- CP-element group 579:  members (6) 
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_sample_completed_
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_update_start_
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/$exit
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Sample/ack
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/$entry
      -- CP-element group 579: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/req
      -- 
    ack_2992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1457_inst_ack_0, ack => concat_CP_34_elements(579)); -- 
    req_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(579), ack => WPIPE_Concat_output_pipe_1457_inst_req_1); -- 
    -- CP-element group 580:  transition  input  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	579 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	581 
    -- CP-element group 580:  members (3) 
      -- CP-element group 580: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_update_completed_
      -- CP-element group 580: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/$exit
      -- CP-element group 580: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1457_Update/ack
      -- 
    ack_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1457_inst_ack_1, ack => concat_CP_34_elements(580)); -- 
    -- CP-element group 581:  join  transition  output  bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	576 
    -- CP-element group 581: 	580 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	582 
    -- CP-element group 581:  members (3) 
      -- CP-element group 581: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_sample_start_
      -- CP-element group 581: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/$entry
      -- CP-element group 581: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/req
      -- 
    req_3005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(581), ack => WPIPE_Concat_output_pipe_1460_inst_req_0); -- 
    concat_cp_element_group_581: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_581"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(576) & concat_CP_34_elements(580);
      gj_concat_cp_element_group_581 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(581), clk => clk, reset => reset); --
    end block;
    -- CP-element group 582:  transition  input  output  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	581 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	583 
    -- CP-element group 582:  members (6) 
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_sample_completed_
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_update_start_
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/$exit
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Sample/ack
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/$entry
      -- CP-element group 582: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/req
      -- 
    ack_3006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 582_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1460_inst_ack_0, ack => concat_CP_34_elements(582)); -- 
    req_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(582), ack => WPIPE_Concat_output_pipe_1460_inst_req_1); -- 
    -- CP-element group 583:  transition  input  bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	582 
    -- CP-element group 583: successors 
    -- CP-element group 583: 	584 
    -- CP-element group 583:  members (3) 
      -- CP-element group 583: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_update_completed_
      -- CP-element group 583: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/$exit
      -- CP-element group 583: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1460_Update/ack
      -- 
    ack_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1460_inst_ack_1, ack => concat_CP_34_elements(583)); -- 
    -- CP-element group 584:  join  transition  output  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	574 
    -- CP-element group 584: 	583 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	585 
    -- CP-element group 584:  members (3) 
      -- CP-element group 584: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/req
      -- 
    req_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(584), ack => WPIPE_Concat_output_pipe_1463_inst_req_0); -- 
    concat_cp_element_group_584: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_584"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(574) & concat_CP_34_elements(583);
      gj_concat_cp_element_group_584 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(584), clk => clk, reset => reset); --
    end block;
    -- CP-element group 585:  transition  input  output  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	584 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	586 
    -- CP-element group 585:  members (6) 
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_sample_completed_
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_update_start_
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/$exit
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Sample/ack
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/$entry
      -- CP-element group 585: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/req
      -- 
    ack_3020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 585_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1463_inst_ack_0, ack => concat_CP_34_elements(585)); -- 
    req_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(585), ack => WPIPE_Concat_output_pipe_1463_inst_req_1); -- 
    -- CP-element group 586:  transition  input  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	585 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	587 
    -- CP-element group 586:  members (3) 
      -- CP-element group 586: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_update_completed_
      -- CP-element group 586: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/$exit
      -- CP-element group 586: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1463_Update/ack
      -- 
    ack_3025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 586_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1463_inst_ack_1, ack => concat_CP_34_elements(586)); -- 
    -- CP-element group 587:  join  transition  output  bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	572 
    -- CP-element group 587: 	586 
    -- CP-element group 587: successors 
    -- CP-element group 587: 	588 
    -- CP-element group 587:  members (3) 
      -- CP-element group 587: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_sample_start_
      -- CP-element group 587: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/$entry
      -- CP-element group 587: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/req
      -- 
    req_3033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(587), ack => WPIPE_Concat_output_pipe_1466_inst_req_0); -- 
    concat_cp_element_group_587: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_587"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(572) & concat_CP_34_elements(586);
      gj_concat_cp_element_group_587 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(587), clk => clk, reset => reset); --
    end block;
    -- CP-element group 588:  transition  input  output  bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	587 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	589 
    -- CP-element group 588:  members (6) 
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_sample_completed_
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_update_start_
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/$exit
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Sample/ack
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/$entry
      -- CP-element group 588: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/req
      -- 
    ack_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1466_inst_ack_0, ack => concat_CP_34_elements(588)); -- 
    req_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(588), ack => WPIPE_Concat_output_pipe_1466_inst_req_1); -- 
    -- CP-element group 589:  transition  input  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	588 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	590 
    -- CP-element group 589:  members (3) 
      -- CP-element group 589: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_update_completed_
      -- CP-element group 589: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/$exit
      -- CP-element group 589: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1466_Update/ack
      -- 
    ack_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 589_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1466_inst_ack_1, ack => concat_CP_34_elements(589)); -- 
    -- CP-element group 590:  join  transition  output  bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	570 
    -- CP-element group 590: 	589 
    -- CP-element group 590: successors 
    -- CP-element group 590: 	591 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_sample_start_
      -- CP-element group 590: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/$entry
      -- CP-element group 590: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/req
      -- 
    req_3047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(590), ack => WPIPE_Concat_output_pipe_1469_inst_req_0); -- 
    concat_cp_element_group_590: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_590"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(570) & concat_CP_34_elements(589);
      gj_concat_cp_element_group_590 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(590), clk => clk, reset => reset); --
    end block;
    -- CP-element group 591:  transition  input  output  bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	590 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	592 
    -- CP-element group 591:  members (6) 
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_sample_completed_
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_update_start_
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/$exit
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Sample/ack
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/$entry
      -- CP-element group 591: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/req
      -- 
    ack_3048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1469_inst_ack_0, ack => concat_CP_34_elements(591)); -- 
    req_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(591), ack => WPIPE_Concat_output_pipe_1469_inst_req_1); -- 
    -- CP-element group 592:  transition  input  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	591 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	593 
    -- CP-element group 592:  members (3) 
      -- CP-element group 592: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_update_completed_
      -- CP-element group 592: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/$exit
      -- CP-element group 592: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1469_Update/ack
      -- 
    ack_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1469_inst_ack_1, ack => concat_CP_34_elements(592)); -- 
    -- CP-element group 593:  join  transition  output  bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	568 
    -- CP-element group 593: 	592 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	594 
    -- CP-element group 593:  members (3) 
      -- CP-element group 593: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_sample_start_
      -- CP-element group 593: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/req
      -- 
    req_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(593), ack => WPIPE_Concat_output_pipe_1472_inst_req_0); -- 
    concat_cp_element_group_593: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_593"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(568) & concat_CP_34_elements(592);
      gj_concat_cp_element_group_593 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(593), clk => clk, reset => reset); --
    end block;
    -- CP-element group 594:  transition  input  output  bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	593 
    -- CP-element group 594: successors 
    -- CP-element group 594: 	595 
    -- CP-element group 594:  members (6) 
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_sample_completed_
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_update_start_
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/$exit
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Sample/ack
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/$entry
      -- CP-element group 594: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/req
      -- 
    ack_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 594_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1472_inst_ack_0, ack => concat_CP_34_elements(594)); -- 
    req_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(594), ack => WPIPE_Concat_output_pipe_1472_inst_req_1); -- 
    -- CP-element group 595:  transition  input  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	594 
    -- CP-element group 595: successors 
    -- CP-element group 595: 	596 
    -- CP-element group 595:  members (3) 
      -- CP-element group 595: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_update_completed_
      -- CP-element group 595: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/$exit
      -- CP-element group 595: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1472_Update/ack
      -- 
    ack_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1472_inst_ack_1, ack => concat_CP_34_elements(595)); -- 
    -- CP-element group 596:  join  transition  output  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	566 
    -- CP-element group 596: 	595 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	597 
    -- CP-element group 596:  members (3) 
      -- CP-element group 596: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_sample_start_
      -- CP-element group 596: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/$entry
      -- CP-element group 596: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/req
      -- 
    req_3075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(596), ack => WPIPE_Concat_output_pipe_1475_inst_req_0); -- 
    concat_cp_element_group_596: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_596"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(566) & concat_CP_34_elements(595);
      gj_concat_cp_element_group_596 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(596), clk => clk, reset => reset); --
    end block;
    -- CP-element group 597:  transition  input  output  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	596 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	598 
    -- CP-element group 597:  members (6) 
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_sample_completed_
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_update_start_
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/$exit
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Sample/ack
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/$entry
      -- CP-element group 597: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/req
      -- 
    ack_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 597_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1475_inst_ack_0, ack => concat_CP_34_elements(597)); -- 
    req_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(597), ack => WPIPE_Concat_output_pipe_1475_inst_req_1); -- 
    -- CP-element group 598:  transition  input  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	597 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	599 
    -- CP-element group 598:  members (3) 
      -- CP-element group 598: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_update_completed_
      -- CP-element group 598: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/$exit
      -- CP-element group 598: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1475_Update/ack
      -- 
    ack_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 598_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1475_inst_ack_1, ack => concat_CP_34_elements(598)); -- 
    -- CP-element group 599:  join  transition  output  bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	564 
    -- CP-element group 599: 	598 
    -- CP-element group 599: successors 
    -- CP-element group 599: 	600 
    -- CP-element group 599:  members (3) 
      -- CP-element group 599: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_sample_start_
      -- CP-element group 599: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/$entry
      -- CP-element group 599: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/req
      -- 
    req_3089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(599), ack => WPIPE_Concat_output_pipe_1478_inst_req_0); -- 
    concat_cp_element_group_599: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_599"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(564) & concat_CP_34_elements(598);
      gj_concat_cp_element_group_599 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(599), clk => clk, reset => reset); --
    end block;
    -- CP-element group 600:  transition  input  output  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	599 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	601 
    -- CP-element group 600:  members (6) 
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_sample_completed_
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_update_start_
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/$exit
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Sample/ack
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/$entry
      -- CP-element group 600: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/req
      -- 
    ack_3090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1478_inst_ack_0, ack => concat_CP_34_elements(600)); -- 
    req_3094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(600), ack => WPIPE_Concat_output_pipe_1478_inst_req_1); -- 
    -- CP-element group 601:  branch  transition  place  input  output  bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	600 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	602 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (17) 
      -- CP-element group 601: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480__exit__
      -- CP-element group 601: 	 branch_block_stmt_23/assign_stmt_1487__entry__
      -- CP-element group 601: 	 branch_block_stmt_23/assign_stmt_1487__exit__
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488__entry__
      -- CP-element group 601: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/$exit
      -- CP-element group 601: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_update_completed_
      -- CP-element group 601: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/$exit
      -- CP-element group 601: 	 branch_block_stmt_23/call_stmt_1372_to_assign_stmt_1480/WPIPE_Concat_output_pipe_1478_Update/ack
      -- CP-element group 601: 	 branch_block_stmt_23/assign_stmt_1487/$entry
      -- CP-element group 601: 	 branch_block_stmt_23/assign_stmt_1487/$exit
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_dead_link/$entry
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_eval_test/$entry
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_eval_test/$exit
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_eval_test/branch_req
      -- CP-element group 601: 	 branch_block_stmt_23/R_cmp381460_1489_place
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_if_link/$entry
      -- CP-element group 601: 	 branch_block_stmt_23/if_stmt_1488_else_link/$entry
      -- 
    ack_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1478_inst_ack_1, ack => concat_CP_34_elements(601)); -- 
    branch_req_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(601), ack => if_stmt_1488_branch_req_0); -- 
    -- CP-element group 602:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	601 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	604 
    -- CP-element group 602: 	605 
    -- CP-element group 602:  members (18) 
      -- CP-element group 602: 	 branch_block_stmt_23/merge_stmt_1494__exit__
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523__entry__
      -- CP-element group 602: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/dummy
      -- CP-element group 602: 	 branch_block_stmt_23/merge_stmt_1494_PhiReqMerge
      -- CP-element group 602: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 602: 	 branch_block_stmt_23/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/whilex_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 602: 	 branch_block_stmt_23/if_stmt_1488_if_link/$exit
      -- CP-element group 602: 	 branch_block_stmt_23/if_stmt_1488_if_link/if_choice_transition
      -- CP-element group 602: 	 branch_block_stmt_23/whilex_xend_bbx_xnph
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_sample_start_
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_update_start_
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/rr
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/cr
      -- 
    if_choice_transition_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 602_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_1, ack => concat_CP_34_elements(602)); -- 
    rr_3128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(602), ack => type_cast_1509_inst_req_0); -- 
    cr_3133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(602), ack => type_cast_1509_inst_req_1); -- 
    -- CP-element group 603:  transition  place  input  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	601 
    -- CP-element group 603: successors 
    -- CP-element group 603: 	674 
    -- CP-element group 603:  members (5) 
      -- CP-element group 603: 	 branch_block_stmt_23/whilex_xend_forx_xend456_PhiReq/$entry
      -- CP-element group 603: 	 branch_block_stmt_23/whilex_xend_forx_xend456_PhiReq/$exit
      -- CP-element group 603: 	 branch_block_stmt_23/if_stmt_1488_else_link/$exit
      -- CP-element group 603: 	 branch_block_stmt_23/if_stmt_1488_else_link/else_choice_transition
      -- CP-element group 603: 	 branch_block_stmt_23/whilex_xend_forx_xend456
      -- 
    else_choice_transition_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_0, ack => concat_CP_34_elements(603)); -- 
    -- CP-element group 604:  transition  input  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	602 
    -- CP-element group 604: successors 
    -- CP-element group 604:  members (3) 
      -- CP-element group 604: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_sample_completed_
      -- CP-element group 604: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/$exit
      -- CP-element group 604: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Sample/ra
      -- 
    ra_3129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_0, ack => concat_CP_34_elements(604)); -- 
    -- CP-element group 605:  transition  place  input  bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	602 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	668 
    -- CP-element group 605:  members (9) 
      -- CP-element group 605: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523__exit__
      -- CP-element group 605: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383
      -- CP-element group 605: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- CP-element group 605: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/$entry
      -- CP-element group 605: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 605: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/$exit
      -- CP-element group 605: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_update_completed_
      -- CP-element group 605: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/$exit
      -- CP-element group 605: 	 branch_block_stmt_23/assign_stmt_1500_to_assign_stmt_1523/type_cast_1509_Update/ca
      -- 
    ca_3134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 605_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_1, ack => concat_CP_34_elements(605)); -- 
    -- CP-element group 606:  transition  input  bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	673 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	651 
    -- CP-element group 606:  members (3) 
      -- CP-element group 606: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_sample_complete
      -- CP-element group 606: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/$exit
      -- CP-element group 606: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/ack
      -- 
    ack_3163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1538_index_offset_ack_0, ack => concat_CP_34_elements(606)); -- 
    -- CP-element group 607:  transition  input  output  bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	673 
    -- CP-element group 607: successors 
    -- CP-element group 607: 	608 
    -- CP-element group 607:  members (11) 
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_sample_start_
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_root_address_calculated
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_offset_calculated
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/$exit
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/ack
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/$entry
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/$exit
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/sum_rename_req
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_base_plus_offset/sum_rename_ack
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/$entry
      -- CP-element group 607: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/req
      -- 
    ack_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1538_index_offset_ack_1, ack => concat_CP_34_elements(607)); -- 
    req_3177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(607), ack => addr_of_1539_final_reg_req_0); -- 
    -- CP-element group 608:  transition  input  bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	607 
    -- CP-element group 608: successors 
    -- CP-element group 608:  members (3) 
      -- CP-element group 608: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_sample_completed_
      -- CP-element group 608: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/$exit
      -- CP-element group 608: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_request/ack
      -- 
    ack_3178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1539_final_reg_ack_0, ack => concat_CP_34_elements(608)); -- 
    -- CP-element group 609:  join  fork  transition  input  output  bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	673 
    -- CP-element group 609: successors 
    -- CP-element group 609: 	610 
    -- CP-element group 609:  members (24) 
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_update_completed_
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/$exit
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/ack
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_sample_start_
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_address_calculated
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_address_calculated
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_root_address_calculated
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_address_resized
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/$exit
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/base_resize_req
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_addr_resize/base_resize_ack
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/$exit
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/sum_rename_req
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_base_plus_offset/sum_rename_ack
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/$exit
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/root_register_req
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_word_addrgen/root_register_ack
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/$entry
      -- CP-element group 609: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/rr
      -- 
    ack_3183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1539_final_reg_ack_1, ack => concat_CP_34_elements(609)); -- 
    rr_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(609), ack => ptr_deref_1543_load_0_req_0); -- 
    -- CP-element group 610:  transition  input  bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	609 
    -- CP-element group 610: successors 
    -- CP-element group 610:  members (5) 
      -- CP-element group 610: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_sample_completed_
      -- CP-element group 610: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/$exit
      -- CP-element group 610: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/$exit
      -- CP-element group 610: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/$exit
      -- CP-element group 610: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Sample/word_access_start/word_0/ra
      -- 
    ra_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 610_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_load_0_ack_0, ack => concat_CP_34_elements(610)); -- 
    -- CP-element group 611:  fork  transition  input  output  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	673 
    -- CP-element group 611: successors 
    -- CP-element group 611: 	612 
    -- CP-element group 611: 	614 
    -- CP-element group 611: 	616 
    -- CP-element group 611: 	618 
    -- CP-element group 611: 	620 
    -- CP-element group 611: 	622 
    -- CP-element group 611: 	624 
    -- CP-element group 611: 	626 
    -- CP-element group 611:  members (33) 
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_update_completed_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/$exit
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/$exit
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/$exit
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/ca
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/$exit
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/merge_req
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/ptr_deref_1543_Merge/merge_ack
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_sample_start_
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/$entry
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/rr
      -- CP-element group 611: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_sample_start_
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 611_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_load_0_ack_1, ack => concat_CP_34_elements(611)); -- 
    rr_3241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1547_inst_req_0); -- 
    rr_3255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1557_inst_req_0); -- 
    rr_3269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1567_inst_req_0); -- 
    rr_3283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1577_inst_req_0); -- 
    rr_3297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1587_inst_req_0); -- 
    rr_3311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1597_inst_req_0); -- 
    rr_3325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1607_inst_req_0); -- 
    rr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(611), ack => type_cast_1617_inst_req_0); -- 
    -- CP-element group 612:  transition  input  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	611 
    -- CP-element group 612: successors 
    -- CP-element group 612:  members (3) 
      -- CP-element group 612: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_sample_completed_
      -- CP-element group 612: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/$exit
      -- CP-element group 612: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Sample/ra
      -- 
    ra_3242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1547_inst_ack_0, ack => concat_CP_34_elements(612)); -- 
    -- CP-element group 613:  transition  input  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	673 
    -- CP-element group 613: successors 
    -- CP-element group 613: 	648 
    -- CP-element group 613:  members (3) 
      -- CP-element group 613: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_update_completed_
      -- CP-element group 613: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/$exit
      -- CP-element group 613: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/ca
      -- 
    ca_3247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 613_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1547_inst_ack_1, ack => concat_CP_34_elements(613)); -- 
    -- CP-element group 614:  transition  input  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	611 
    -- CP-element group 614: successors 
    -- CP-element group 614:  members (3) 
      -- CP-element group 614: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_sample_completed_
      -- CP-element group 614: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/$exit
      -- CP-element group 614: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Sample/ra
      -- 
    ra_3256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 614_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_0, ack => concat_CP_34_elements(614)); -- 
    -- CP-element group 615:  transition  input  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	673 
    -- CP-element group 615: successors 
    -- CP-element group 615: 	645 
    -- CP-element group 615:  members (3) 
      -- CP-element group 615: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_update_completed_
      -- CP-element group 615: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/$exit
      -- CP-element group 615: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/ca
      -- 
    ca_3261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_1, ack => concat_CP_34_elements(615)); -- 
    -- CP-element group 616:  transition  input  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	611 
    -- CP-element group 616: successors 
    -- CP-element group 616:  members (3) 
      -- CP-element group 616: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_sample_completed_
      -- CP-element group 616: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/$exit
      -- CP-element group 616: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Sample/ra
      -- 
    ra_3270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_0, ack => concat_CP_34_elements(616)); -- 
    -- CP-element group 617:  transition  input  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	673 
    -- CP-element group 617: successors 
    -- CP-element group 617: 	642 
    -- CP-element group 617:  members (3) 
      -- CP-element group 617: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_update_completed_
      -- CP-element group 617: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/$exit
      -- CP-element group 617: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/ca
      -- 
    ca_3275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_1, ack => concat_CP_34_elements(617)); -- 
    -- CP-element group 618:  transition  input  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	611 
    -- CP-element group 618: successors 
    -- CP-element group 618:  members (3) 
      -- CP-element group 618: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_sample_completed_
      -- CP-element group 618: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/$exit
      -- CP-element group 618: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Sample/ra
      -- 
    ra_3284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_0, ack => concat_CP_34_elements(618)); -- 
    -- CP-element group 619:  transition  input  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	673 
    -- CP-element group 619: successors 
    -- CP-element group 619: 	639 
    -- CP-element group 619:  members (3) 
      -- CP-element group 619: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_update_completed_
      -- CP-element group 619: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/$exit
      -- CP-element group 619: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/ca
      -- 
    ca_3289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 619_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_1, ack => concat_CP_34_elements(619)); -- 
    -- CP-element group 620:  transition  input  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	611 
    -- CP-element group 620: successors 
    -- CP-element group 620:  members (3) 
      -- CP-element group 620: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_sample_completed_
      -- CP-element group 620: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/$exit
      -- CP-element group 620: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Sample/ra
      -- 
    ra_3298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_0, ack => concat_CP_34_elements(620)); -- 
    -- CP-element group 621:  transition  input  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	673 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	636 
    -- CP-element group 621:  members (3) 
      -- CP-element group 621: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_update_completed_
      -- CP-element group 621: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/$exit
      -- CP-element group 621: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/ca
      -- 
    ca_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_1, ack => concat_CP_34_elements(621)); -- 
    -- CP-element group 622:  transition  input  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	611 
    -- CP-element group 622: successors 
    -- CP-element group 622:  members (3) 
      -- CP-element group 622: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/ra
      -- CP-element group 622: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Sample/$exit
      -- CP-element group 622: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_sample_completed_
      -- 
    ra_3312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_0, ack => concat_CP_34_elements(622)); -- 
    -- CP-element group 623:  transition  input  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	673 
    -- CP-element group 623: successors 
    -- CP-element group 623: 	633 
    -- CP-element group 623:  members (3) 
      -- CP-element group 623: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/ca
      -- CP-element group 623: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/$exit
      -- CP-element group 623: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_update_completed_
      -- 
    ca_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1597_inst_ack_1, ack => concat_CP_34_elements(623)); -- 
    -- CP-element group 624:  transition  input  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	611 
    -- CP-element group 624: successors 
    -- CP-element group 624:  members (3) 
      -- CP-element group 624: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_sample_completed_
      -- CP-element group 624: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/$exit
      -- CP-element group 624: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Sample/ra
      -- 
    ra_3326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_0, ack => concat_CP_34_elements(624)); -- 
    -- CP-element group 625:  transition  input  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	673 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	630 
    -- CP-element group 625:  members (3) 
      -- CP-element group 625: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_update_completed_
      -- CP-element group 625: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/$exit
      -- CP-element group 625: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/ca
      -- 
    ca_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1607_inst_ack_1, ack => concat_CP_34_elements(625)); -- 
    -- CP-element group 626:  transition  input  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	611 
    -- CP-element group 626: successors 
    -- CP-element group 626:  members (3) 
      -- CP-element group 626: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_sample_completed_
      -- CP-element group 626: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/ra
      -- CP-element group 626: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Sample/$exit
      -- 
    ra_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_0, ack => concat_CP_34_elements(626)); -- 
    -- CP-element group 627:  transition  input  output  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	673 
    -- CP-element group 627: successors 
    -- CP-element group 627: 	628 
    -- CP-element group 627:  members (6) 
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_sample_start_
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/ca
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/$exit
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_update_completed_
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/$entry
      -- CP-element group 627: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/req
      -- 
    ca_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_1, ack => concat_CP_34_elements(627)); -- 
    req_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(627), ack => WPIPE_Concat_output_pipe_1619_inst_req_0); -- 
    -- CP-element group 628:  transition  input  output  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	627 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	629 
    -- CP-element group 628:  members (6) 
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_sample_completed_
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_update_start_
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/req
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/$entry
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/ack
      -- CP-element group 628: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Sample/$exit
      -- 
    ack_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1619_inst_ack_0, ack => concat_CP_34_elements(628)); -- 
    req_3358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(628), ack => WPIPE_Concat_output_pipe_1619_inst_req_1); -- 
    -- CP-element group 629:  transition  input  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	628 
    -- CP-element group 629: successors 
    -- CP-element group 629: 	630 
    -- CP-element group 629:  members (3) 
      -- CP-element group 629: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_update_completed_
      -- CP-element group 629: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/ack
      -- CP-element group 629: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1619_Update/$exit
      -- 
    ack_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1619_inst_ack_1, ack => concat_CP_34_elements(629)); -- 
    -- CP-element group 630:  join  transition  output  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	625 
    -- CP-element group 630: 	629 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	631 
    -- CP-element group 630:  members (3) 
      -- CP-element group 630: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/req
      -- CP-element group 630: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/$entry
      -- CP-element group 630: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_sample_start_
      -- 
    req_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(630), ack => WPIPE_Concat_output_pipe_1622_inst_req_0); -- 
    concat_cp_element_group_630: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_630"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(625) & concat_CP_34_elements(629);
      gj_concat_cp_element_group_630 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(630), clk => clk, reset => reset); --
    end block;
    -- CP-element group 631:  transition  input  output  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	630 
    -- CP-element group 631: successors 
    -- CP-element group 631: 	632 
    -- CP-element group 631:  members (6) 
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/req
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/$entry
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/ack
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Sample/$exit
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_update_start_
      -- CP-element group 631: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_sample_completed_
      -- 
    ack_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1622_inst_ack_0, ack => concat_CP_34_elements(631)); -- 
    req_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(631), ack => WPIPE_Concat_output_pipe_1622_inst_req_1); -- 
    -- CP-element group 632:  transition  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	631 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	633 
    -- CP-element group 632:  members (3) 
      -- CP-element group 632: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/ack
      -- CP-element group 632: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_Update/$exit
      -- CP-element group 632: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1622_update_completed_
      -- 
    ack_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1622_inst_ack_1, ack => concat_CP_34_elements(632)); -- 
    -- CP-element group 633:  join  transition  output  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	623 
    -- CP-element group 633: 	632 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	634 
    -- CP-element group 633:  members (3) 
      -- CP-element group 633: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/req
      -- CP-element group 633: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/$entry
      -- CP-element group 633: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_sample_start_
      -- 
    req_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(633), ack => WPIPE_Concat_output_pipe_1625_inst_req_0); -- 
    concat_cp_element_group_633: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_633"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(623) & concat_CP_34_elements(632);
      gj_concat_cp_element_group_633 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(633), clk => clk, reset => reset); --
    end block;
    -- CP-element group 634:  transition  input  output  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	633 
    -- CP-element group 634: successors 
    -- CP-element group 634: 	635 
    -- CP-element group 634:  members (6) 
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/req
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/ack
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Sample/$exit
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_update_start_
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/$entry
      -- CP-element group 634: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_sample_completed_
      -- 
    ack_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 634_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1625_inst_ack_0, ack => concat_CP_34_elements(634)); -- 
    req_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(634), ack => WPIPE_Concat_output_pipe_1625_inst_req_1); -- 
    -- CP-element group 635:  transition  input  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	634 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	636 
    -- CP-element group 635:  members (3) 
      -- CP-element group 635: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/ack
      -- CP-element group 635: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_Update/$exit
      -- CP-element group 635: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1625_update_completed_
      -- 
    ack_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1625_inst_ack_1, ack => concat_CP_34_elements(635)); -- 
    -- CP-element group 636:  join  transition  output  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	621 
    -- CP-element group 636: 	635 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	637 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_sample_start_
      -- CP-element group 636: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/$entry
      -- CP-element group 636: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/req
      -- 
    req_3395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(636), ack => WPIPE_Concat_output_pipe_1628_inst_req_0); -- 
    concat_cp_element_group_636: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_636"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(621) & concat_CP_34_elements(635);
      gj_concat_cp_element_group_636 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(636), clk => clk, reset => reset); --
    end block;
    -- CP-element group 637:  transition  input  output  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	636 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	638 
    -- CP-element group 637:  members (6) 
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/req
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/$entry
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/ack
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_sample_completed_
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_update_start_
      -- CP-element group 637: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Sample/$exit
      -- 
    ack_3396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1628_inst_ack_0, ack => concat_CP_34_elements(637)); -- 
    req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(637), ack => WPIPE_Concat_output_pipe_1628_inst_req_1); -- 
    -- CP-element group 638:  transition  input  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	637 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	639 
    -- CP-element group 638:  members (3) 
      -- CP-element group 638: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/$exit
      -- CP-element group 638: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_update_completed_
      -- CP-element group 638: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1628_Update/ack
      -- 
    ack_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 638_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1628_inst_ack_1, ack => concat_CP_34_elements(638)); -- 
    -- CP-element group 639:  join  transition  output  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	619 
    -- CP-element group 639: 	638 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	640 
    -- CP-element group 639:  members (3) 
      -- CP-element group 639: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/req
      -- CP-element group 639: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/$entry
      -- CP-element group 639: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_sample_start_
      -- 
    req_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(639), ack => WPIPE_Concat_output_pipe_1631_inst_req_0); -- 
    concat_cp_element_group_639: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_639"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(619) & concat_CP_34_elements(638);
      gj_concat_cp_element_group_639 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(639), clk => clk, reset => reset); --
    end block;
    -- CP-element group 640:  transition  input  output  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	639 
    -- CP-element group 640: successors 
    -- CP-element group 640: 	641 
    -- CP-element group 640:  members (6) 
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/ack
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/$entry
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Sample/$exit
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/req
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_sample_completed_
      -- CP-element group 640: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_update_start_
      -- 
    ack_3410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1631_inst_ack_0, ack => concat_CP_34_elements(640)); -- 
    req_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(640), ack => WPIPE_Concat_output_pipe_1631_inst_req_1); -- 
    -- CP-element group 641:  transition  input  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	640 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	642 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/$exit
      -- CP-element group 641: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_update_completed_
      -- CP-element group 641: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1631_Update/ack
      -- 
    ack_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 641_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1631_inst_ack_1, ack => concat_CP_34_elements(641)); -- 
    -- CP-element group 642:  join  transition  output  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	617 
    -- CP-element group 642: 	641 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	643 
    -- CP-element group 642:  members (3) 
      -- CP-element group 642: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/req
      -- CP-element group 642: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/$entry
      -- CP-element group 642: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_sample_start_
      -- 
    req_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(642), ack => WPIPE_Concat_output_pipe_1634_inst_req_0); -- 
    concat_cp_element_group_642: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_642"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(617) & concat_CP_34_elements(641);
      gj_concat_cp_element_group_642 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(642), clk => clk, reset => reset); --
    end block;
    -- CP-element group 643:  transition  input  output  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	642 
    -- CP-element group 643: successors 
    -- CP-element group 643: 	644 
    -- CP-element group 643:  members (6) 
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/req
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/$entry
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/ack
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Sample/$exit
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_update_start_
      -- CP-element group 643: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_sample_completed_
      -- 
    ack_3424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1634_inst_ack_0, ack => concat_CP_34_elements(643)); -- 
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(643), ack => WPIPE_Concat_output_pipe_1634_inst_req_1); -- 
    -- CP-element group 644:  transition  input  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	643 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644:  members (3) 
      -- CP-element group 644: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/ack
      -- CP-element group 644: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_Update/$exit
      -- CP-element group 644: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1634_update_completed_
      -- 
    ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 644_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1634_inst_ack_1, ack => concat_CP_34_elements(644)); -- 
    -- CP-element group 645:  join  transition  output  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	615 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	646 
    -- CP-element group 645:  members (3) 
      -- CP-element group 645: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/req
      -- CP-element group 645: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/$entry
      -- CP-element group 645: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_sample_start_
      -- 
    req_3437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(645), ack => WPIPE_Concat_output_pipe_1637_inst_req_0); -- 
    concat_cp_element_group_645: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_645"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(615) & concat_CP_34_elements(644);
      gj_concat_cp_element_group_645 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(645), clk => clk, reset => reset); --
    end block;
    -- CP-element group 646:  transition  input  output  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	645 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646:  members (6) 
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/req
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/$entry
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/ack
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Sample/$exit
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_update_start_
      -- CP-element group 646: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_sample_completed_
      -- 
    ack_3438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1637_inst_ack_0, ack => concat_CP_34_elements(646)); -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(646), ack => WPIPE_Concat_output_pipe_1637_inst_req_1); -- 
    -- CP-element group 647:  transition  input  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	648 
    -- CP-element group 647:  members (3) 
      -- CP-element group 647: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/ack
      -- CP-element group 647: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_Update/$exit
      -- CP-element group 647: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1637_update_completed_
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1637_inst_ack_1, ack => concat_CP_34_elements(647)); -- 
    -- CP-element group 648:  join  transition  output  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	613 
    -- CP-element group 648: 	647 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (3) 
      -- CP-element group 648: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/req
      -- CP-element group 648: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/$entry
      -- CP-element group 648: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_sample_start_
      -- 
    req_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(648), ack => WPIPE_Concat_output_pipe_1640_inst_req_0); -- 
    concat_cp_element_group_648: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_648"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(613) & concat_CP_34_elements(647);
      gj_concat_cp_element_group_648 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(648), clk => clk, reset => reset); --
    end block;
    -- CP-element group 649:  transition  input  output  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649: 	650 
    -- CP-element group 649:  members (6) 
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/req
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/$exit
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Sample/ack
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/$entry
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_update_start_
      -- CP-element group 649: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_sample_completed_
      -- 
    ack_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1640_inst_ack_0, ack => concat_CP_34_elements(649)); -- 
    req_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(649), ack => WPIPE_Concat_output_pipe_1640_inst_req_1); -- 
    -- CP-element group 650:  transition  input  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	649 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	651 
    -- CP-element group 650:  members (3) 
      -- CP-element group 650: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/$exit
      -- CP-element group 650: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_Update/ack
      -- CP-element group 650: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/WPIPE_Concat_output_pipe_1640_update_completed_
      -- 
    ack_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 650_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1640_inst_ack_1, ack => concat_CP_34_elements(650)); -- 
    -- CP-element group 651:  branch  join  transition  place  output  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	606 
    -- CP-element group 651: 	650 
    -- CP-element group 651: successors 
    -- CP-element group 651: 	652 
    -- CP-element group 651: 	653 
    -- CP-element group 651:  members (10) 
      -- CP-element group 651: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653__exit__
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654__entry__
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_else_link/$entry
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_if_link/$entry
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_eval_test/branch_req
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_dead_link/$entry
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_eval_test/$entry
      -- CP-element group 651: 	 branch_block_stmt_23/if_stmt_1654_eval_test/$exit
      -- CP-element group 651: 	 branch_block_stmt_23/R_exitcond1_1655_place
      -- CP-element group 651: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/$exit
      -- 
    branch_req_3465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(651), ack => if_stmt_1654_branch_req_0); -- 
    concat_cp_element_group_651: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_651"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(606) & concat_CP_34_elements(650);
      gj_concat_cp_element_group_651 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(651), clk => clk, reset => reset); --
    end block;
    -- CP-element group 652:  merge  transition  place  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	651 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	674 
    -- CP-element group 652:  members (13) 
      -- CP-element group 652: 	 branch_block_stmt_23/merge_stmt_1660__exit__
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456
      -- CP-element group 652: 	 branch_block_stmt_23/if_stmt_1654_if_link/if_choice_transition
      -- CP-element group 652: 	 branch_block_stmt_23/merge_stmt_1660_PhiReqMerge
      -- CP-element group 652: 	 branch_block_stmt_23/if_stmt_1654_if_link/$exit
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456_PhiReq/$exit
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xend456x_xloopexit_forx_xend456_PhiReq/$entry
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit
      -- CP-element group 652: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/dummy
      -- CP-element group 652: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/$exit
      -- CP-element group 652: 	 branch_block_stmt_23/merge_stmt_1660_PhiAck/$entry
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit_PhiReq/$exit
      -- CP-element group 652: 	 branch_block_stmt_23/forx_xbody383_forx_xend456x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_3470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1654_branch_ack_1, ack => concat_CP_34_elements(652)); -- 
    -- CP-element group 653:  fork  transition  place  input  output  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	651 
    -- CP-element group 653: successors 
    -- CP-element group 653: 	669 
    -- CP-element group 653: 	670 
    -- CP-element group 653:  members (12) 
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/if_stmt_1654_else_link/$exit
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383
      -- CP-element group 653: 	 branch_block_stmt_23/if_stmt_1654_else_link/else_choice_transition
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/cr
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/rr
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/$entry
      -- CP-element group 653: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/$entry
      -- 
    else_choice_transition_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 653_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1654_branch_ack_0, ack => concat_CP_34_elements(653)); -- 
    cr_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(653), ack => type_cast_1532_inst_req_1); -- 
    rr_3691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(653), ack => type_cast_1532_inst_req_0); -- 
    -- CP-element group 654:  merge  branch  transition  place  output  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	76 
    -- CP-element group 654: 	121 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	77 
    -- CP-element group 654: 	78 
    -- CP-element group 654:  members (17) 
      -- CP-element group 654: 	 branch_block_stmt_23/merge_stmt_316__exit__
      -- CP-element group 654: 	 branch_block_stmt_23/assign_stmt_322__entry__
      -- CP-element group 654: 	 branch_block_stmt_23/assign_stmt_322__exit__
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323__entry__
      -- CP-element group 654: 	 branch_block_stmt_23/assign_stmt_322/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/assign_stmt_322/$exit
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_dead_link/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_eval_test/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_eval_test/$exit
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_eval_test/branch_req
      -- CP-element group 654: 	 branch_block_stmt_23/R_cmp175463_324_place
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_if_link/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/if_stmt_323_else_link/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/merge_stmt_316_PhiAck/$exit
      -- CP-element group 654: 	 branch_block_stmt_23/merge_stmt_316_PhiAck/$entry
      -- CP-element group 654: 	 branch_block_stmt_23/merge_stmt_316_PhiReqMerge
      -- CP-element group 654: 	 branch_block_stmt_23/merge_stmt_316_PhiAck/dummy
      -- 
    branch_req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(654), ack => if_stmt_323_branch_req_0); -- 
    concat_CP_34_elements(654) <= OrReduce(concat_CP_34_elements(76) & concat_CP_34_elements(121));
    -- CP-element group 655:  transition  output  delay-element  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	80 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	659 
    -- CP-element group 655:  members (5) 
      -- CP-element group 655: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_req
      -- CP-element group 655: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_381_konst_delay_trans
      -- CP-element group 655: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/$exit
      -- CP-element group 655: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_377/$exit
      -- CP-element group 655: 	 branch_block_stmt_23/bbx_xnph469_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_377_req_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_377_req_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(655), ack => phi_stmt_377_req_0); -- 
    -- Element group concat_CP_34_elements(655) is a control-delay.
    cp_element_655_delay: control_delay_element  generic map(name => " 655_delay", delay_value => 1)  port map(req => concat_CP_34_elements(80), ack => concat_CP_34_elements(655), clk => clk, reset =>reset);
    -- CP-element group 656:  transition  input  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	122 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	658 
    -- CP-element group 656:  members (2) 
      -- CP-element group 656: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Sample/ra
      -- CP-element group 656: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Sample/$exit
      -- 
    ra_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_0, ack => concat_CP_34_elements(656)); -- 
    -- CP-element group 657:  transition  input  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	122 
    -- CP-element group 657: successors 
    -- CP-element group 657: 	658 
    -- CP-element group 657:  members (2) 
      -- CP-element group 657: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Update/ca
      -- CP-element group 657: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/Update/$exit
      -- 
    ca_3547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 657_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_1, ack => concat_CP_34_elements(657)); -- 
    -- CP-element group 658:  join  transition  output  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	656 
    -- CP-element group 658: 	657 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (6) 
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_req
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/SplitProtocol/$exit
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/type_cast_383/$exit
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/phi_stmt_377_sources/$exit
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_377/$exit
      -- CP-element group 658: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_377_req_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_377_req_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(658), ack => phi_stmt_377_req_1); -- 
    concat_cp_element_group_658: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_658"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(656) & concat_CP_34_elements(657);
      gj_concat_cp_element_group_658 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(658), clk => clk, reset => reset); --
    end block;
    -- CP-element group 659:  merge  transition  place  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	655 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	660 
    -- CP-element group 659:  members (2) 
      -- CP-element group 659: 	 branch_block_stmt_23/merge_stmt_376_PhiReqMerge
      -- CP-element group 659: 	 branch_block_stmt_23/merge_stmt_376_PhiAck/$entry
      -- 
    concat_CP_34_elements(659) <= OrReduce(concat_CP_34_elements(655) & concat_CP_34_elements(658));
    -- CP-element group 660:  fork  transition  place  input  output  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	659 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	81 
    -- CP-element group 660: 	82 
    -- CP-element group 660: 	84 
    -- CP-element group 660: 	85 
    -- CP-element group 660: 	88 
    -- CP-element group 660: 	92 
    -- CP-element group 660: 	96 
    -- CP-element group 660: 	100 
    -- CP-element group 660: 	104 
    -- CP-element group 660: 	108 
    -- CP-element group 660: 	112 
    -- CP-element group 660: 	116 
    -- CP-element group 660: 	119 
    -- CP-element group 660:  members (56) 
      -- CP-element group 660: 	 branch_block_stmt_23/merge_stmt_376__exit__
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539__entry__
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/word_0/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/word_0/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/word_access_complete/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_410_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_resized_1
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_scaled_1
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_computed_1
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_resize_1/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_resize_1/$exit
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_resize_1/index_resize_req
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_resize_1/index_resize_ack
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_scale_1/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_scale_1/$exit
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_scale_1/scale_rename_req
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_index_scale_1/scale_rename_ack
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_update_start
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Sample/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Sample/req
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/array_obj_ref_389_final_index_sum_regn_Update/req
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_complete/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/addr_of_390_complete/req
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_sample_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Sample/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/RPIPE_Concat_input_pipe_393_Sample/rr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_397_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_428_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_446_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_464_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_482_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_500_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/type_cast_518_Update/cr
      -- CP-element group 660: 	 branch_block_stmt_23/assign_stmt_391_to_assign_stmt_539/ptr_deref_526_update_start_
      -- CP-element group 660: 	 branch_block_stmt_23/merge_stmt_376_PhiAck/phi_stmt_377_ack
      -- CP-element group 660: 	 branch_block_stmt_23/merge_stmt_376_PhiAck/$exit
      -- 
    phi_stmt_377_ack_3553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_377_ack_0, ack => concat_CP_34_elements(660)); -- 
    cr_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => ptr_deref_526_store_0_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_410_inst_req_1); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => array_obj_ref_389_index_offset_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => array_obj_ref_389_index_offset_req_1); -- 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => addr_of_390_final_reg_req_1); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => RPIPE_Concat_input_pipe_393_inst_req_0); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_397_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_428_inst_req_1); -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_446_inst_req_1); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_464_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_482_inst_req_1); -- 
    cr_922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_500_inst_req_1); -- 
    cr_950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(660), ack => type_cast_518_inst_req_1); -- 
    -- CP-element group 661:  transition  output  delay-element  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	124 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	665 
    -- CP-element group 661:  members (5) 
      -- CP-element group 661: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_598_konst_delay_trans
      -- CP-element group 661: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_req
      -- CP-element group 661: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/$exit
      -- CP-element group 661: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_594/$exit
      -- CP-element group 661: 	 branch_block_stmt_23/bbx_xnph465_forx_xbody177_PhiReq/$exit
      -- 
    phi_stmt_594_req_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_594_req_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(661), ack => phi_stmt_594_req_0); -- 
    -- Element group concat_CP_34_elements(661) is a control-delay.
    cp_element_661_delay: control_delay_element  generic map(name => " 661_delay", delay_value => 1)  port map(req => concat_CP_34_elements(124), ack => concat_CP_34_elements(661), clk => clk, reset =>reset);
    -- CP-element group 662:  transition  input  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	166 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	664 
    -- CP-element group 662:  members (2) 
      -- CP-element group 662: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Sample/$exit
      -- CP-element group 662: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Sample/ra
      -- 
    ra_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 662_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_600_inst_ack_0, ack => concat_CP_34_elements(662)); -- 
    -- CP-element group 663:  transition  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	166 
    -- CP-element group 663: successors 
    -- CP-element group 663: 	664 
    -- CP-element group 663:  members (2) 
      -- CP-element group 663: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Update/ca
      -- CP-element group 663: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/Update/$exit
      -- 
    ca_3601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_600_inst_ack_1, ack => concat_CP_34_elements(663)); -- 
    -- CP-element group 664:  join  transition  output  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	662 
    -- CP-element group 664: 	663 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	665 
    -- CP-element group 664:  members (6) 
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_sources/type_cast_600/SplitProtocol/$exit
      -- CP-element group 664: 	 branch_block_stmt_23/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_594/phi_stmt_594_req
      -- 
    phi_stmt_594_req_3602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_594_req_3602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(664), ack => phi_stmt_594_req_1); -- 
    concat_cp_element_group_664: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_664"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(662) & concat_CP_34_elements(663);
      gj_concat_cp_element_group_664 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(664), clk => clk, reset => reset); --
    end block;
    -- CP-element group 665:  merge  transition  place  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	661 
    -- CP-element group 665: 	664 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	666 
    -- CP-element group 665:  members (2) 
      -- CP-element group 665: 	 branch_block_stmt_23/merge_stmt_593_PhiReqMerge
      -- CP-element group 665: 	 branch_block_stmt_23/merge_stmt_593_PhiAck/$entry
      -- 
    concat_CP_34_elements(665) <= OrReduce(concat_CP_34_elements(661) & concat_CP_34_elements(664));
    -- CP-element group 666:  fork  transition  place  input  output  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	665 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	125 
    -- CP-element group 666: 	126 
    -- CP-element group 666: 	128 
    -- CP-element group 666: 	129 
    -- CP-element group 666: 	132 
    -- CP-element group 666: 	136 
    -- CP-element group 666: 	140 
    -- CP-element group 666: 	144 
    -- CP-element group 666: 	148 
    -- CP-element group 666: 	152 
    -- CP-element group 666: 	156 
    -- CP-element group 666: 	160 
    -- CP-element group 666: 	163 
    -- CP-element group 666:  members (56) 
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_computed_1
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_scaled_1
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/word_0/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/word_0/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_resized_1
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_sample_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/merge_stmt_593__exit__
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756__entry__
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_scale_1/scale_rename_ack
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_scale_1/scale_rename_req
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_scale_1/$exit
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_scale_1/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_resize_1/index_resize_ack
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_resize_1/index_resize_req
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/word_access_complete/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_627_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/ptr_deref_743_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_complete/req
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/addr_of_607_complete/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_645_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_663_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_735_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Sample/rr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_resize_1/$exit
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/RPIPE_Concat_input_pipe_610_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_index_resize_1/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_699_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_681_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Update/cr
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_614_update_start_
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/type_cast_717_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Update/req
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Update/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Sample/req
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_Sample/$entry
      -- CP-element group 666: 	 branch_block_stmt_23/assign_stmt_608_to_assign_stmt_756/array_obj_ref_606_final_index_sum_regn_update_start
      -- CP-element group 666: 	 branch_block_stmt_23/merge_stmt_593_PhiAck/phi_stmt_594_ack
      -- CP-element group 666: 	 branch_block_stmt_23/merge_stmt_593_PhiAck/$exit
      -- 
    phi_stmt_594_ack_3607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_594_ack_0, ack => concat_CP_34_elements(666)); -- 
    cr_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => ptr_deref_743_store_0_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_627_inst_req_1); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_645_inst_req_1); -- 
    req_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => addr_of_607_final_reg_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_663_inst_req_1); -- 
    cr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_699_inst_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_681_inst_req_1); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_614_inst_req_1); -- 
    cr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_735_inst_req_1); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => RPIPE_Concat_input_pipe_610_inst_req_0); -- 
    cr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => type_cast_717_inst_req_1); -- 
    req_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => array_obj_ref_606_index_offset_req_1); -- 
    req_1065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(666), ack => array_obj_ref_606_index_offset_req_0); -- 
    -- CP-element group 667:  merge  fork  transition  place  output  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	78 
    -- CP-element group 667: 	165 
    -- CP-element group 667: successors 
    -- CP-element group 667: 	167 
    -- CP-element group 667: 	168 
    -- CP-element group 667:  members (13) 
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_update_start_
      -- CP-element group 667: 	 branch_block_stmt_23/merge_stmt_765__exit__
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768__entry__
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/$entry
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/ccr
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Update/$entry
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/crr
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_Sample/$entry
      -- CP-element group 667: 	 branch_block_stmt_23/call_stmt_768/call_stmt_768_sample_start_
      -- CP-element group 667: 	 branch_block_stmt_23/merge_stmt_765_PhiReqMerge
      -- CP-element group 667: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/dummy
      -- CP-element group 667: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/$exit
      -- CP-element group 667: 	 branch_block_stmt_23/merge_stmt_765_PhiAck/$entry
      -- 
    ccr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(667), ack => call_stmt_768_call_req_1); -- 
    crr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(667), ack => call_stmt_768_call_req_0); -- 
    concat_CP_34_elements(667) <= OrReduce(concat_CP_34_elements(78) & concat_CP_34_elements(165));
    -- CP-element group 668:  transition  output  delay-element  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	605 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	672 
    -- CP-element group 668:  members (5) 
      -- CP-element group 668: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 668: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/$exit
      -- CP-element group 668: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/$exit
      -- CP-element group 668: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1530_konst_delay_trans
      -- CP-element group 668: 	 branch_block_stmt_23/bbx_xnph_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- 
    phi_stmt_1526_req_3672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_3672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(668), ack => phi_stmt_1526_req_0); -- 
    -- Element group concat_CP_34_elements(668) is a control-delay.
    cp_element_668_delay: control_delay_element  generic map(name => " 668_delay", delay_value => 1)  port map(req => concat_CP_34_elements(605), ack => concat_CP_34_elements(668), clk => clk, reset =>reset);
    -- CP-element group 669:  transition  input  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	653 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	671 
    -- CP-element group 669:  members (2) 
      -- CP-element group 669: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/ra
      -- CP-element group 669: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Sample/$exit
      -- 
    ra_3692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1532_inst_ack_0, ack => concat_CP_34_elements(669)); -- 
    -- CP-element group 670:  transition  input  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	653 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	671 
    -- CP-element group 670:  members (2) 
      -- CP-element group 670: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/ca
      -- CP-element group 670: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/Update/$exit
      -- 
    ca_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 670_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1532_inst_ack_1, ack => concat_CP_34_elements(670)); -- 
    -- CP-element group 671:  join  transition  output  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	669 
    -- CP-element group 671: 	670 
    -- CP-element group 671: successors 
    -- CP-element group 671: 	672 
    -- CP-element group 671:  members (6) 
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/$exit
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/$exit
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532/SplitProtocol/$exit
      -- CP-element group 671: 	 branch_block_stmt_23/forx_xbody383_forx_xbody383_PhiReq/$exit
      -- 
    phi_stmt_1526_req_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(671), ack => phi_stmt_1526_req_1); -- 
    concat_cp_element_group_671: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_671"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_34_elements(669) & concat_CP_34_elements(670);
      gj_concat_cp_element_group_671 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_34_elements(671), clk => clk, reset => reset); --
    end block;
    -- CP-element group 672:  merge  transition  place  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	668 
    -- CP-element group 672: 	671 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	673 
    -- CP-element group 672:  members (2) 
      -- CP-element group 672: 	 branch_block_stmt_23/merge_stmt_1525_PhiReqMerge
      -- CP-element group 672: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/$entry
      -- 
    concat_CP_34_elements(672) <= OrReduce(concat_CP_34_elements(668) & concat_CP_34_elements(671));
    -- CP-element group 673:  fork  transition  place  input  output  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	672 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	606 
    -- CP-element group 673: 	607 
    -- CP-element group 673: 	609 
    -- CP-element group 673: 	611 
    -- CP-element group 673: 	613 
    -- CP-element group 673: 	615 
    -- CP-element group 673: 	617 
    -- CP-element group 673: 	619 
    -- CP-element group 673: 	621 
    -- CP-element group 673: 	623 
    -- CP-element group 673: 	625 
    -- CP-element group 673: 	627 
    -- CP-element group 673:  members (53) 
      -- CP-element group 673: 	 branch_block_stmt_23/merge_stmt_1525__exit__
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653__entry__
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1607_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1617_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/phi_stmt_1526_ack
      -- CP-element group 673: 	 branch_block_stmt_23/merge_stmt_1525_PhiAck/$exit
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resized_1
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scaled_1
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_computed_1
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/$exit
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/index_resize_req
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_resize_1/index_resize_ack
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/$exit
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/scale_rename_req
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_index_scale_1/scale_rename_ack
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_update_start
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Sample/req
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/array_obj_ref_1538_final_index_sum_regn_Update/req
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/addr_of_1539_complete/req
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/ptr_deref_1543_Update/word_access_complete/word_0/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1547_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1557_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1567_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1577_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_update_start_
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/$entry
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1587_Update/cr
      -- CP-element group 673: 	 branch_block_stmt_23/assign_stmt_1540_to_assign_stmt_1653/type_cast_1597_update_start_
      -- 
    phi_stmt_1526_ack_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 673_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1526_ack_0, ack => concat_CP_34_elements(673)); -- 
    cr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1617_inst_req_1); -- 
    cr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1607_inst_req_1); -- 
    cr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1597_inst_req_1); -- 
    req_3162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => array_obj_ref_1538_index_offset_req_0); -- 
    req_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => array_obj_ref_1538_index_offset_req_1); -- 
    req_3182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => addr_of_1539_final_reg_req_1); -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => ptr_deref_1543_load_0_req_1); -- 
    cr_3246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1547_inst_req_1); -- 
    cr_3260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1557_inst_req_1); -- 
    cr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1567_inst_req_1); -- 
    cr_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1577_inst_req_1); -- 
    cr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_34_elements(673), ack => type_cast_1587_inst_req_1); -- 
    -- CP-element group 674:  merge  transition  place  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	603 
    -- CP-element group 674: 	652 
    -- CP-element group 674: successors 
    -- CP-element group 674:  members (16) 
      -- CP-element group 674: 	 $exit
      -- CP-element group 674: 	 branch_block_stmt_23/$exit
      -- CP-element group 674: 	 branch_block_stmt_23/branch_block_stmt_23__exit__
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1662__exit__
      -- CP-element group 674: 	 branch_block_stmt_23/return__
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1664__exit__
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1662_PhiReqMerge
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1664_PhiReqMerge
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/dummy
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/$entry
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/$exit
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1662_PhiAck/dummy
      -- CP-element group 674: 	 branch_block_stmt_23/return___PhiReq/$entry
      -- CP-element group 674: 	 branch_block_stmt_23/return___PhiReq/$exit
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/$exit
      -- CP-element group 674: 	 branch_block_stmt_23/merge_stmt_1664_PhiAck/$entry
      -- 
    concat_CP_34_elements(674) <= OrReduce(concat_CP_34_elements(603) & concat_CP_34_elements(652));
    concat_do_while_stmt_817_terminator_2805: loop_terminator -- 
      generic map (name => " concat_do_while_stmt_817_terminator_2805", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_CP_34_elements(173),loop_continue => concat_CP_34_elements(553),loop_terminate => concat_CP_34_elements(552),loop_back => concat_CP_34_elements(171),loop_exit => concat_CP_34_elements(170),clk => clk, reset => reset); -- 
    phi_stmt_819_phi_seq_1463_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(186);
      concat_CP_34_elements(191)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(195);
      concat_CP_34_elements(192)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(196);
      concat_CP_34_elements(187) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(188);
      concat_CP_34_elements(197)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(197);
      concat_CP_34_elements(198)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(199);
      concat_CP_34_elements(189) <= phi_mux_reqs(1);
      phi_stmt_819_phi_seq_1463 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_819_phi_seq_1463") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(178), 
          phi_sample_ack => concat_CP_34_elements(184), 
          phi_update_req => concat_CP_34_elements(180), 
          phi_update_ack => concat_CP_34_elements(185), 
          phi_mux_ack => concat_CP_34_elements(190), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_824_phi_seq_1507_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(207);
      concat_CP_34_elements(212)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(216);
      concat_CP_34_elements(213)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(217);
      concat_CP_34_elements(208) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(209);
      concat_CP_34_elements(218)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(218);
      concat_CP_34_elements(219)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(220);
      concat_CP_34_elements(210) <= phi_mux_reqs(1);
      phi_stmt_824_phi_seq_1507 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_824_phi_seq_1507") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(203), 
          phi_sample_ack => concat_CP_34_elements(204), 
          phi_update_req => concat_CP_34_elements(205), 
          phi_update_ack => concat_CP_34_elements(206), 
          phi_mux_ack => concat_CP_34_elements(211), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_829_phi_seq_1551_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(228);
      concat_CP_34_elements(233)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(237);
      concat_CP_34_elements(234)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(238);
      concat_CP_34_elements(229) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(230);
      concat_CP_34_elements(239)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(239);
      concat_CP_34_elements(240)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(241);
      concat_CP_34_elements(231) <= phi_mux_reqs(1);
      phi_stmt_829_phi_seq_1551 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_829_phi_seq_1551") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(224), 
          phi_sample_ack => concat_CP_34_elements(225), 
          phi_update_req => concat_CP_34_elements(226), 
          phi_update_ack => concat_CP_34_elements(227), 
          phi_mux_ack => concat_CP_34_elements(232), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_834_phi_seq_1595_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(249);
      concat_CP_34_elements(254)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(258);
      concat_CP_34_elements(255)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(259);
      concat_CP_34_elements(250) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(251);
      concat_CP_34_elements(260)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(260);
      concat_CP_34_elements(261)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(262);
      concat_CP_34_elements(252) <= phi_mux_reqs(1);
      phi_stmt_834_phi_seq_1595 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_834_phi_seq_1595") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(245), 
          phi_sample_ack => concat_CP_34_elements(246), 
          phi_update_req => concat_CP_34_elements(247), 
          phi_update_ack => concat_CP_34_elements(248), 
          phi_mux_ack => concat_CP_34_elements(253), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_839_phi_seq_1639_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_CP_34_elements(270);
      concat_CP_34_elements(275)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_CP_34_elements(279);
      concat_CP_34_elements(276)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_CP_34_elements(280);
      concat_CP_34_elements(271) <= phi_mux_reqs(0);
      triggers(1)  <= concat_CP_34_elements(272);
      concat_CP_34_elements(281)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_CP_34_elements(281);
      concat_CP_34_elements(282)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_CP_34_elements(283);
      concat_CP_34_elements(273) <= phi_mux_reqs(1);
      phi_stmt_839_phi_seq_1639 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_839_phi_seq_1639") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_CP_34_elements(266), 
          phi_sample_ack => concat_CP_34_elements(267), 
          phi_update_req => concat_CP_34_elements(268), 
          phi_update_ack => concat_CP_34_elements(269), 
          phi_mux_ack => concat_CP_34_elements(274), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1415_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_CP_34_elements(174);
        preds(1)  <= concat_CP_34_elements(175);
        entry_tmerge_1415 : transition_merge -- 
          generic map(name => " entry_tmerge_1415")
          port map (preds => preds, symbol_out => concat_CP_34_elements(176));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1152_1152_delayed_2_0_1254 : std_logic_vector(15 downto 0);
    signal MUX_1166_wire : std_logic_vector(15 downto 0);
    signal MUX_1168_1168_delayed_2_0_1282 : std_logic_vector(15 downto 0);
    signal MUX_1181_wire : std_logic_vector(15 downto 0);
    signal MUX_1185_1185_delayed_2_0_1306 : std_logic_vector(15 downto 0);
    signal MUX_1196_wire : std_logic_vector(15 downto 0);
    signal MUX_1202_1202_delayed_2_0_1332 : std_logic_vector(15 downto 0);
    signal MUX_1261_wire : std_logic_vector(15 downto 0);
    signal MUX_1289_wire : std_logic_vector(15 downto 0);
    signal MUX_1315_wire : std_logic_vector(15 downto 0);
    signal MUX_1341_wire : std_logic_vector(15 downto 0);
    signal MUX_963_wire : std_logic_vector(15 downto 0);
    signal MUX_978_wire : std_logic_vector(15 downto 0);
    signal MUX_993_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1024_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1061_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1227_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1358_wire : std_logic_vector(0 downto 0);
    signal R_idxprom247_875_resized : std_logic_vector(13 downto 0);
    signal R_idxprom247_875_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom251_898_resized : std_logic_vector(13 downto 0);
    signal R_idxprom251_898_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom273_1078_resized : std_logic_vector(13 downto 0);
    signal R_idxprom273_1078_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom277_1101_resized : std_logic_vector(13 downto 0);
    signal R_idxprom277_1101_scaled : std_logic_vector(13 downto 0);
    signal R_indvar476_605_resized : std_logic_vector(13 downto 0);
    signal R_indvar476_605_scaled : std_logic_vector(13 downto 0);
    signal R_indvar489_388_resized : std_logic_vector(13 downto 0);
    signal R_indvar489_388_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1537_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1537_scaled : std_logic_vector(13 downto 0);
    signal add12_74 : std_logic_vector(31 downto 0);
    signal add131_416 : std_logic_vector(63 downto 0);
    signal add137_434 : std_logic_vector(63 downto 0);
    signal add143_452 : std_logic_vector(63 downto 0);
    signal add149_470 : std_logic_vector(63 downto 0);
    signal add155_488 : std_logic_vector(63 downto 0);
    signal add161_506 : std_logic_vector(63 downto 0);
    signal add167_524 : std_logic_vector(63 downto 0);
    signal add187_633 : std_logic_vector(63 downto 0);
    signal add193_651 : std_logic_vector(63 downto 0);
    signal add199_669 : std_logic_vector(63 downto 0);
    signal add205_687 : std_logic_vector(63 downto 0);
    signal add211_705 : std_logic_vector(63 downto 0);
    signal add217_723 : std_logic_vector(63 downto 0);
    signal add21_99 : std_logic_vector(31 downto 0);
    signal add223_741 : std_logic_vector(63 downto 0);
    signal add30_124 : std_logic_vector(31 downto 0);
    signal add39_149 : std_logic_vector(31 downto 0);
    signal add48_174 : std_logic_vector(31 downto 0);
    signal add57_199 : std_logic_vector(31 downto 0);
    signal add66_224 : std_logic_vector(31 downto 0);
    signal add75_249 : std_logic_vector(31 downto 0);
    signal add_49 : std_logic_vector(31 downto 0);
    signal add_inp1x_x0_980 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_824 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_866_delayed_1_0_866 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_907_delayed_1_0_925 : std_logic_vector(15 downto 0);
    signal add_inp1x_x1_at_entry_796 : std_logic_vector(15 downto 0);
    signal add_inp2x_x0506_1263 : std_logic_vector(15 downto 0);
    signal add_inp2x_x0x_xph_1183 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_1015_delayed_3_0_1069 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_1056_delayed_3_0_1128 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_829 : std_logic_vector(15 downto 0);
    signal add_inp2x_x1_at_entry_801 : std_logic_vector(15 downto 0);
    signal add_outx_x0_1032_delayed_2_0_1092 : std_logic_vector(15 downto 0);
    signal add_outx_x0_1063_delayed_2_0_1138 : std_logic_vector(15 downto 0);
    signal add_outx_x0_965 : std_logic_vector(15 downto 0);
    signal add_outx_x1_819 : std_logic_vector(15 downto 0);
    signal add_outx_x1_883_delayed_1_0_889 : std_logic_vector(15 downto 0);
    signal add_outx_x1_914_delayed_1_0_935 : std_logic_vector(15 downto 0);
    signal add_outx_x1_at_entry_790 : std_logic_vector(15 downto 0);
    signal add_outx_x2504_1291 : std_logic_vector(15 downto 0);
    signal add_outx_x2x_xph_1168 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1079_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1102_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1538_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_389_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_606_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_899_root_address : std_logic_vector(13 downto 0);
    signal arrayidx227_608 : std_logic_vector(31 downto 0);
    signal arrayidx248_878 : std_logic_vector(31 downto 0);
    signal arrayidx252_894_delayed_6_0_907 : std_logic_vector(31 downto 0);
    signal arrayidx252_901 : std_logic_vector(31 downto 0);
    signal arrayidx274_1081 : std_logic_vector(31 downto 0);
    signal arrayidx278_1043_delayed_6_0_1110 : std_logic_vector(31 downto 0);
    signal arrayidx278_1104 : std_logic_vector(31 downto 0);
    signal arrayidx388_1540 : std_logic_vector(31 downto 0);
    signal arrayidx_391 : std_logic_vector(31 downto 0);
    signal call10_65 : std_logic_vector(7 downto 0);
    signal call124_394 : std_logic_vector(7 downto 0);
    signal call128_407 : std_logic_vector(7 downto 0);
    signal call134_425 : std_logic_vector(7 downto 0);
    signal call140_443 : std_logic_vector(7 downto 0);
    signal call146_461 : std_logic_vector(7 downto 0);
    signal call14_77 : std_logic_vector(7 downto 0);
    signal call152_479 : std_logic_vector(7 downto 0);
    signal call158_497 : std_logic_vector(7 downto 0);
    signal call164_515 : std_logic_vector(7 downto 0);
    signal call180_611 : std_logic_vector(7 downto 0);
    signal call184_624 : std_logic_vector(7 downto 0);
    signal call190_642 : std_logic_vector(7 downto 0);
    signal call196_660 : std_logic_vector(7 downto 0);
    signal call19_90 : std_logic_vector(7 downto 0);
    signal call202_678 : std_logic_vector(7 downto 0);
    signal call208_696 : std_logic_vector(7 downto 0);
    signal call214_714 : std_logic_vector(7 downto 0);
    signal call220_732 : std_logic_vector(7 downto 0);
    signal call233_768 : std_logic_vector(63 downto 0);
    signal call23_102 : std_logic_vector(7 downto 0);
    signal call28_115 : std_logic_vector(7 downto 0);
    signal call2_40 : std_logic_vector(7 downto 0);
    signal call310_1372 : std_logic_vector(63 downto 0);
    signal call32_127 : std_logic_vector(7 downto 0);
    signal call37_140 : std_logic_vector(7 downto 0);
    signal call41_152 : std_logic_vector(7 downto 0);
    signal call46_165 : std_logic_vector(7 downto 0);
    signal call50_177 : std_logic_vector(7 downto 0);
    signal call55_190 : std_logic_vector(7 downto 0);
    signal call59_202 : std_logic_vector(7 downto 0);
    signal call5_52 : std_logic_vector(7 downto 0);
    signal call64_215 : std_logic_vector(7 downto 0);
    signal call68_227 : std_logic_vector(7 downto 0);
    signal call73_240 : std_logic_vector(7 downto 0);
    signal call_26 : std_logic_vector(7 downto 0);
    signal cmp175463_322 : std_logic_vector(0 downto 0);
    signal cmp244_853 : std_logic_vector(0 downto 0);
    signal cmp263_1009 : std_logic_vector(0 downto 0);
    signal cmp269_1046 : std_logic_vector(0 downto 0);
    signal cmp297_1212 : std_logic_vector(0 downto 0);
    signal cmp305_1352 : std_logic_vector(0 downto 0);
    signal cmp381460_1487 : std_logic_vector(0 downto 0);
    signal cmp467_307 : std_logic_vector(0 downto 0);
    signal conv11_69 : std_logic_vector(31 downto 0);
    signal conv125_398 : std_logic_vector(63 downto 0);
    signal conv130_411 : std_logic_vector(63 downto 0);
    signal conv136_429 : std_logic_vector(63 downto 0);
    signal conv142_447 : std_logic_vector(63 downto 0);
    signal conv148_465 : std_logic_vector(63 downto 0);
    signal conv154_483 : std_logic_vector(63 downto 0);
    signal conv160_501 : std_logic_vector(63 downto 0);
    signal conv166_519 : std_logic_vector(63 downto 0);
    signal conv17_81 : std_logic_vector(31 downto 0);
    signal conv181_615 : std_logic_vector(63 downto 0);
    signal conv186_628 : std_logic_vector(63 downto 0);
    signal conv192_646 : std_logic_vector(63 downto 0);
    signal conv198_664 : std_logic_vector(63 downto 0);
    signal conv1_31 : std_logic_vector(31 downto 0);
    signal conv204_682 : std_logic_vector(63 downto 0);
    signal conv20_94 : std_logic_vector(31 downto 0);
    signal conv210_700 : std_logic_vector(63 downto 0);
    signal conv216_718 : std_logic_vector(63 downto 0);
    signal conv222_736 : std_logic_vector(63 downto 0);
    signal conv234_1369 : std_logic_vector(63 downto 0);
    signal conv241_848 : std_logic_vector(31 downto 0);
    signal conv243_775 : std_logic_vector(31 downto 0);
    signal conv260_1000 : std_logic_vector(31 downto 0);
    signal conv266_1037 : std_logic_vector(31 downto 0);
    signal conv268_781 : std_logic_vector(31 downto 0);
    signal conv26_106 : std_logic_vector(31 downto 0);
    signal conv294_1203 : std_logic_vector(31 downto 0);
    signal conv29_119 : std_logic_vector(31 downto 0);
    signal conv302_1347 : std_logic_vector(31 downto 0);
    signal conv311_1377 : std_logic_vector(63 downto 0);
    signal conv317_1386 : std_logic_vector(7 downto 0);
    signal conv323_1396 : std_logic_vector(7 downto 0);
    signal conv329_1406 : std_logic_vector(7 downto 0);
    signal conv335_1416 : std_logic_vector(7 downto 0);
    signal conv341_1426 : std_logic_vector(7 downto 0);
    signal conv347_1436 : std_logic_vector(7 downto 0);
    signal conv353_1446 : std_logic_vector(7 downto 0);
    signal conv359_1456 : std_logic_vector(7 downto 0);
    signal conv35_131 : std_logic_vector(31 downto 0);
    signal conv38_144 : std_logic_vector(31 downto 0);
    signal conv393_1548 : std_logic_vector(7 downto 0);
    signal conv399_1558 : std_logic_vector(7 downto 0);
    signal conv3_44 : std_logic_vector(31 downto 0);
    signal conv405_1568 : std_logic_vector(7 downto 0);
    signal conv411_1578 : std_logic_vector(7 downto 0);
    signal conv417_1588 : std_logic_vector(7 downto 0);
    signal conv423_1598 : std_logic_vector(7 downto 0);
    signal conv429_1608 : std_logic_vector(7 downto 0);
    signal conv435_1618 : std_logic_vector(7 downto 0);
    signal conv44_156 : std_logic_vector(31 downto 0);
    signal conv47_169 : std_logic_vector(31 downto 0);
    signal conv53_181 : std_logic_vector(31 downto 0);
    signal conv56_194 : std_logic_vector(31 downto 0);
    signal conv62_206 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv71_231 : std_logic_vector(31 downto 0);
    signal conv74_244 : std_logic_vector(31 downto 0);
    signal conv8_56 : std_logic_vector(31 downto 0);
    signal count_inp1x_x0_995 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_834 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_900_delayed_1_0_915 : std_logic_vector(15 downto 0);
    signal count_inp1x_x1_at_entry_806 : std_logic_vector(15 downto 0);
    signal count_inp1x_x2_1317 : std_logic_vector(15 downto 0);
    signal count_inp2x_x0x_xph_1198 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_1049_delayed_3_0_1118 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_839 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_990_delayed_2_0_1032 : std_logic_vector(15 downto 0);
    signal count_inp2x_x1_at_entry_811 : std_logic_vector(15 downto 0);
    signal count_inp2x_x2_1343 : std_logic_vector(15 downto 0);
    signal exitcond1_1653 : std_logic_vector(0 downto 0);
    signal exitcond2_539 : std_logic_vector(0 downto 0);
    signal exitcond_756 : std_logic_vector(0 downto 0);
    signal iNsTr_19_361 : std_logic_vector(63 downto 0);
    signal iNsTr_32_578 : std_logic_vector(63 downto 0);
    signal iNsTr_79_1510 : std_logic_vector(63 downto 0);
    signal idxprom247_871 : std_logic_vector(63 downto 0);
    signal idxprom251_894 : std_logic_vector(63 downto 0);
    signal idxprom273_1074 : std_logic_vector(63 downto 0);
    signal idxprom277_1097 : std_logic_vector(63 downto 0);
    signal ifx_xend300_whilex_xend_taken_1355 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_950 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_968_delayed_1_0_1003 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_975_delayed_1_0_1012 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_980_delayed_1_0_1020 : std_logic_vector(0 downto 0);
    signal ifx_xend_ifx_xend300_taken_1026 : std_logic_vector(0 downto 0);
    signal ifx_xend_landx_xlhsx_xtrue_taken_1017 : std_logic_vector(0 downto 0);
    signal ifx_xthen271_exec_guard_1025_delayed_7_0_1084 : std_logic_vector(0 downto 0);
    signal ifx_xthen271_exec_guard_1042_delayed_13_0_1107 : std_logic_vector(0 downto 0);
    signal ifx_xthen271_exec_guard_1066 : std_logic_vector(0 downto 0);
    signal ifx_xthen271_landx_xlhsx_xtrue292_taken_1148 : std_logic_vector(0 downto 0);
    signal ifx_xthen299_exec_guard_1232 : std_logic_vector(0 downto 0);
    signal ifx_xthen299_ifx_xend300_taken_1235 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_863 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_876_delayed_7_0_881 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_893_delayed_13_0_904 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend_taken_945 : std_logic_vector(0 downto 0);
    signal inc254_922 : std_logic_vector(15 downto 0);
    signal inc256_932 : std_logic_vector(15 downto 0);
    signal inc258_942 : std_logic_vector(15 downto 0);
    signal inc280_1125 : std_logic_vector(15 downto 0);
    signal inc282_1135 : std_logic_vector(15 downto 0);
    signal inc284_1145 : std_logic_vector(15 downto 0);
    signal indvar476_594 : std_logic_vector(63 downto 0);
    signal indvar489_377 : std_logic_vector(63 downto 0);
    signal indvar_1526 : std_logic_vector(63 downto 0);
    signal indvarx_xnext477_751 : std_logic_vector(63 downto 0);
    signal indvarx_xnext490_534 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1648 : std_logic_vector(63 downto 0);
    signal landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1206 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1215 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1223 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue292_exec_guard_1153 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue292_ifx_xend300_taken_1229 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue292_ifx_xthen299_taken_1220 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_1029 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1040 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_ifx_xthen271_taken_1054 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063 : std_logic_vector(0 downto 0);
    signal mul100_274 : std_logic_vector(31 downto 0);
    signal mul103_279 : std_logic_vector(31 downto 0);
    signal mul109_284 : std_logic_vector(31 downto 0);
    signal mul116_295 : std_logic_vector(31 downto 0);
    signal mul85_259 : std_logic_vector(31 downto 0);
    signal mul91_264 : std_logic_vector(31 downto 0);
    signal mul94_269 : std_logic_vector(31 downto 0);
    signal mul_254 : std_logic_vector(31 downto 0);
    signal ptr_deref_1088_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1088_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1088_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1113_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1113_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1113_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1543_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1543_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_526_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_526_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_526_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_526_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_526_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_526_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_743_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_743_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_743_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_743_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_743_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_743_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_885_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_885_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_885_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_885_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_885_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_910_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_910_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_910_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_910_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_910_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_910_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl127_404 : std_logic_vector(63 downto 0);
    signal shl133_422 : std_logic_vector(63 downto 0);
    signal shl139_440 : std_logic_vector(63 downto 0);
    signal shl145_458 : std_logic_vector(63 downto 0);
    signal shl151_476 : std_logic_vector(63 downto 0);
    signal shl157_494 : std_logic_vector(63 downto 0);
    signal shl163_512 : std_logic_vector(63 downto 0);
    signal shl183_621 : std_logic_vector(63 downto 0);
    signal shl189_639 : std_logic_vector(63 downto 0);
    signal shl18_87 : std_logic_vector(31 downto 0);
    signal shl195_657 : std_logic_vector(63 downto 0);
    signal shl201_675 : std_logic_vector(63 downto 0);
    signal shl207_693 : std_logic_vector(63 downto 0);
    signal shl213_711 : std_logic_vector(63 downto 0);
    signal shl219_729 : std_logic_vector(63 downto 0);
    signal shl27_112 : std_logic_vector(31 downto 0);
    signal shl36_137 : std_logic_vector(31 downto 0);
    signal shl45_162 : std_logic_vector(31 downto 0);
    signal shl54_187 : std_logic_vector(31 downto 0);
    signal shl63_212 : std_logic_vector(31 downto 0);
    signal shl72_237 : std_logic_vector(31 downto 0);
    signal shl9_62 : std_logic_vector(31 downto 0);
    signal shl_37 : std_logic_vector(31 downto 0);
    signal shr117458_301 : std_logic_vector(31 downto 0);
    signal shr304_787 : std_logic_vector(31 downto 0);
    signal shr320_1392 : std_logic_vector(63 downto 0);
    signal shr326_1402 : std_logic_vector(63 downto 0);
    signal shr332_1412 : std_logic_vector(63 downto 0);
    signal shr338_1422 : std_logic_vector(63 downto 0);
    signal shr344_1432 : std_logic_vector(63 downto 0);
    signal shr350_1442 : std_logic_vector(63 downto 0);
    signal shr356_1452 : std_logic_vector(63 downto 0);
    signal shr396_1554 : std_logic_vector(63 downto 0);
    signal shr402_1564 : std_logic_vector(63 downto 0);
    signal shr408_1574 : std_logic_vector(63 downto 0);
    signal shr414_1584 : std_logic_vector(63 downto 0);
    signal shr420_1594 : std_logic_vector(63 downto 0);
    signal shr426_1604 : std_logic_vector(63 downto 0);
    signal shr432_1614 : std_logic_vector(63 downto 0);
    signal shr457_290 : std_logic_vector(31 downto 0);
    signal sub_1382 : std_logic_vector(63 downto 0);
    signal tmp249_886 : std_logic_vector(63 downto 0);
    signal tmp275_1089 : std_logic_vector(63 downto 0);
    signal tmp389_1544 : std_logic_vector(63 downto 0);
    signal tmp471x_xop_1506 : std_logic_vector(31 downto 0);
    signal tmp472_1500 : std_logic_vector(0 downto 0);
    signal tmp475_1523 : std_logic_vector(63 downto 0);
    signal tmp479_551 : std_logic_vector(31 downto 0);
    signal tmp481_556 : std_logic_vector(31 downto 0);
    signal tmp482_562 : std_logic_vector(31 downto 0);
    signal tmp482x_xop_574 : std_logic_vector(31 downto 0);
    signal tmp483_568 : std_logic_vector(0 downto 0);
    signal tmp487_591 : std_logic_vector(63 downto 0);
    signal tmp492_334 : std_logic_vector(31 downto 0);
    signal tmp494_339 : std_logic_vector(31 downto 0);
    signal tmp495_345 : std_logic_vector(31 downto 0);
    signal tmp495x_xop_357 : std_logic_vector(31 downto 0);
    signal tmp496_351 : std_logic_vector(0 downto 0);
    signal tmp500_374 : std_logic_vector(63 downto 0);
    signal type_cast_1082_1082_delayed_2_0_1157 : std_logic_vector(15 downto 0);
    signal type_cast_1094_1094_delayed_3_0_1172 : std_logic_vector(15 downto 0);
    signal type_cast_1106_1106_delayed_3_0_1187 : std_logic_vector(15 downto 0);
    signal type_cast_110_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1143_1143_delayed_1_0_1239 : std_logic_vector(15 downto 0);
    signal type_cast_1143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1146_1146_delayed_1_0_1243 : std_logic_vector(15 downto 0);
    signal type_cast_1149_1149_delayed_2_0_1247 : std_logic_vector(15 downto 0);
    signal type_cast_1159_1159_delayed_1_0_1267 : std_logic_vector(15 downto 0);
    signal type_cast_1161_wire : std_logic_vector(15 downto 0);
    signal type_cast_1162_1162_delayed_1_0_1271 : std_logic_vector(15 downto 0);
    signal type_cast_1165_1165_delayed_1_0_1275 : std_logic_vector(15 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1176_wire : std_logic_vector(15 downto 0);
    signal type_cast_1179_1179_delayed_3_0_1295 : std_logic_vector(15 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1182_1182_delayed_1_0_1299 : std_logic_vector(15 downto 0);
    signal type_cast_1191_wire : std_logic_vector(15 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1196_1196_delayed_1_0_1321 : std_logic_vector(15 downto 0);
    signal type_cast_1199_1199_delayed_2_0_1325 : std_logic_vector(15 downto 0);
    signal type_cast_1252_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1280_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1304_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1337_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_135_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1367_wire : std_logic_vector(63 downto 0);
    signal type_cast_1375_wire : std_logic_vector(63 downto 0);
    signal type_cast_1390_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1410_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1498_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1504_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1514_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1521_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1532_wire : std_logic_vector(63 downto 0);
    signal type_cast_1552_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1572_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1592_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1602_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1646_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_235_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_288_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_299_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_305_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_343_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_349_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_355_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_35_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_365_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_372_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_383_wire : std_logic_vector(63 downto 0);
    signal type_cast_402_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_438_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_492_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_510_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_560_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_572_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_598_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_600_wire : std_logic_vector(63 downto 0);
    signal type_cast_60_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_619_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_637_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_655_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_673_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_691_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_709_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_727_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_749_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_779_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_785_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_822_wire : std_logic_vector(15 downto 0);
    signal type_cast_827_wire : std_logic_vector(15 downto 0);
    signal type_cast_832_wire : std_logic_vector(15 downto 0);
    signal type_cast_837_wire : std_logic_vector(15 downto 0);
    signal type_cast_842_wire : std_logic_vector(15 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_930_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_933_933_delayed_1_0_954 : std_logic_vector(15 downto 0);
    signal type_cast_940_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_945_945_delayed_1_0_969 : std_logic_vector(15 downto 0);
    signal type_cast_957_957_delayed_1_0_984 : std_logic_vector(15 downto 0);
    signal type_cast_958_wire : std_logic_vector(15 downto 0);
    signal type_cast_962_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_973_wire : std_logic_vector(15 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_988_wire : std_logic_vector(15 downto 0);
    signal type_cast_992_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_ifx_xend_taken_860 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xthen_taken_856 : std_logic_vector(0 downto 0);
    signal xx_xop502_584 : std_logic_vector(63 downto 0);
    signal xx_xop503_367 : std_logic_vector(63 downto 0);
    signal xx_xop_1516 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    add_inp1x_x1_at_entry_796 <= "0000000000000000";
    add_inp2x_x1_at_entry_801 <= "0000000000000000";
    add_outx_x1_at_entry_790 <= "0000000000000000";
    array_obj_ref_1079_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1079_resized_base_address <= "00000000000000";
    array_obj_ref_1102_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1102_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1102_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1102_resized_base_address <= "00000000000000";
    array_obj_ref_1538_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1538_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1538_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1538_resized_base_address <= "00000000000000";
    array_obj_ref_389_constant_part_of_offset <= "00000000000000";
    array_obj_ref_389_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_389_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_389_resized_base_address <= "00000000000000";
    array_obj_ref_606_constant_part_of_offset <= "00000000000000";
    array_obj_ref_606_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_606_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_606_resized_base_address <= "00000000000000";
    array_obj_ref_876_constant_part_of_offset <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_876_resized_base_address <= "00000000000000";
    array_obj_ref_899_constant_part_of_offset <= "00000000000000";
    array_obj_ref_899_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_899_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_899_resized_base_address <= "00000000000000";
    count_inp1x_x1_at_entry_806 <= "0000000000000000";
    count_inp2x_x1_at_entry_811 <= "0000000000000000";
    ptr_deref_1088_word_offset_0 <= "00000000000000";
    ptr_deref_1113_word_offset_0 <= "00000000000000";
    ptr_deref_1543_word_offset_0 <= "00000000000000";
    ptr_deref_526_word_offset_0 <= "00000000000000";
    ptr_deref_743_word_offset_0 <= "00000000000000";
    ptr_deref_885_word_offset_0 <= "00000000000000";
    ptr_deref_910_word_offset_0 <= "00000000000000";
    type_cast_110_wire_constant <= "00000000000000000000000000001000";
    type_cast_1123_wire_constant <= "0000000000000001";
    type_cast_1133_wire_constant <= "0000000000000001";
    type_cast_1143_wire_constant <= "0000000000000001";
    type_cast_1165_wire_constant <= "0000000000000000";
    type_cast_1180_wire_constant <= "0000000000000000";
    type_cast_1195_wire_constant <= "0000000000000000";
    type_cast_1252_wire_constant <= "0000000000000000";
    type_cast_1280_wire_constant <= "0000000000000000";
    type_cast_1304_wire_constant <= "0000000000000000";
    type_cast_1311_wire_constant <= "0000000000000000";
    type_cast_1330_wire_constant <= "0000000000000000";
    type_cast_1337_wire_constant <= "0000000000000000";
    type_cast_135_wire_constant <= "00000000000000000000000000001000";
    type_cast_1390_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1400_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1430_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1485_wire_constant <= "00000000000000000000000000000111";
    type_cast_1498_wire_constant <= "00000000000000000000000000000001";
    type_cast_1504_wire_constant <= "11111111111111111111111111111111";
    type_cast_1514_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1521_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1552_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1562_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1572_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1592_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1602_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_160_wire_constant <= "00000000000000000000000000001000";
    type_cast_1612_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1646_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_185_wire_constant <= "00000000000000000000000000001000";
    type_cast_210_wire_constant <= "00000000000000000000000000001000";
    type_cast_235_wire_constant <= "00000000000000000000000000001000";
    type_cast_288_wire_constant <= "00000000000000000000000000000011";
    type_cast_299_wire_constant <= "00000000000000000000000000000011";
    type_cast_305_wire_constant <= "00000000000000000000000000000111";
    type_cast_320_wire_constant <= "00000000000000000000000000000111";
    type_cast_343_wire_constant <= "00000000000000000000000000000011";
    type_cast_349_wire_constant <= "00000000000000000000000000000001";
    type_cast_355_wire_constant <= "11111111111111111111111111111111";
    type_cast_35_wire_constant <= "00000000000000000000000000001000";
    type_cast_365_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_381_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_402_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_456_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_474_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_492_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_510_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_560_wire_constant <= "00000000000000000000000000000011";
    type_cast_566_wire_constant <= "00000000000000000000000000000001";
    type_cast_572_wire_constant <= "11111111111111111111111111111111";
    type_cast_582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_598_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_60_wire_constant <= "00000000000000000000000000001000";
    type_cast_619_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_637_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_655_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_673_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_691_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_709_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_727_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_749_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_773_wire_constant <= "00000000000000001111111111111111";
    type_cast_779_wire_constant <= "00000000000000001111111111111111";
    type_cast_785_wire_constant <= "00000000000000000000000000000011";
    type_cast_85_wire_constant <= "00000000000000000000000000001000";
    type_cast_920_wire_constant <= "0000000000000001";
    type_cast_930_wire_constant <= "0000000000000001";
    type_cast_940_wire_constant <= "0000000000000001";
    type_cast_962_wire_constant <= "0000000000000000";
    type_cast_977_wire_constant <= "0000000000000000";
    type_cast_992_wire_constant <= "0000000000000000";
    phi_stmt_1526: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1530_wire_constant & type_cast_1532_wire;
      req <= phi_stmt_1526_req_0 & phi_stmt_1526_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1526",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1526_ack_0,
          idata => idata,
          odata => indvar_1526,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1526
    phi_stmt_377: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_381_wire_constant & type_cast_383_wire;
      req <= phi_stmt_377_req_0 & phi_stmt_377_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_377",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_377_ack_0,
          idata => idata,
          odata => indvar489_377,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_377
    phi_stmt_594: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_598_wire_constant & type_cast_600_wire;
      req <= phi_stmt_594_req_0 & phi_stmt_594_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_594",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_594_ack_0,
          idata => idata,
          odata => indvar476_594,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_594
    phi_stmt_819: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_822_wire & add_outx_x1_at_entry_790;
      req <= phi_stmt_819_req_0 & phi_stmt_819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_819",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_819_ack_0,
          idata => idata,
          odata => add_outx_x1_819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_819
    phi_stmt_824: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_827_wire & add_inp1x_x1_at_entry_796;
      req <= phi_stmt_824_req_0 & phi_stmt_824_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_824",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_824_ack_0,
          idata => idata,
          odata => add_inp1x_x1_824,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_824
    phi_stmt_829: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_832_wire & add_inp2x_x1_at_entry_801;
      req <= phi_stmt_829_req_0 & phi_stmt_829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_829",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_829_ack_0,
          idata => idata,
          odata => add_inp2x_x1_829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_829
    phi_stmt_834: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_837_wire & count_inp1x_x1_at_entry_806;
      req <= phi_stmt_834_req_0 & phi_stmt_834_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_834",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_834_ack_0,
          idata => idata,
          odata => count_inp1x_x1_834,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_834
    phi_stmt_839: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_842_wire & count_inp2x_x1_at_entry_811;
      req <= phi_stmt_839_req_0 & phi_stmt_839_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_839",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_839_ack_0,
          idata => idata,
          odata => count_inp2x_x1_839,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_839
    -- flow-through select operator MUX_1166_inst
    MUX_1166_wire <= type_cast_1082_1082_delayed_2_0_1157 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063(0) /=  '0') else type_cast_1165_wire_constant;
    -- flow-through select operator MUX_1167_inst
    add_outx_x2x_xph_1168 <= type_cast_1161_wire when (ifx_xthen271_landx_xlhsx_xtrue292_taken_1148(0) /=  '0') else MUX_1166_wire;
    -- flow-through select operator MUX_1181_inst
    MUX_1181_wire <= type_cast_1094_1094_delayed_3_0_1172 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063(0) /=  '0') else type_cast_1180_wire_constant;
    -- flow-through select operator MUX_1182_inst
    add_inp2x_x0x_xph_1183 <= type_cast_1176_wire when (ifx_xthen271_landx_xlhsx_xtrue292_taken_1148(0) /=  '0') else MUX_1181_wire;
    -- flow-through select operator MUX_1196_inst
    MUX_1196_wire <= type_cast_1106_1106_delayed_3_0_1187 when (landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063(0) /=  '0') else type_cast_1195_wire_constant;
    -- flow-through select operator MUX_1197_inst
    count_inp2x_x0x_xph_1198 <= type_cast_1191_wire when (ifx_xthen271_landx_xlhsx_xtrue292_taken_1148(0) /=  '0') else MUX_1196_wire;
    MUX_1253_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1253_inst_req_0;
      MUX_1253_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1253_inst_req_1;
      MUX_1253_inst_ack_1<= update_ack(0);
      MUX_1253_inst: SelectSplitProtocol generic map(name => "MUX_1253_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1149_1149_delayed_2_0_1247, y => type_cast_1252_wire_constant, sel => ifx_xend_ifx_xend300_taken_1026, z => MUX_1152_1152_delayed_2_0_1254, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1261_inst
    MUX_1261_wire <= type_cast_1146_1146_delayed_1_0_1243 when (landx_xlhsx_xtrue292_ifx_xend300_taken_1229(0) /=  '0') else MUX_1152_1152_delayed_2_0_1254;
    -- flow-through select operator MUX_1262_inst
    add_inp2x_x0506_1263 <= type_cast_1143_1143_delayed_1_0_1239 when (ifx_xthen299_ifx_xend300_taken_1235(0) /=  '0') else MUX_1261_wire;
    MUX_1281_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1281_inst_req_0;
      MUX_1281_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1281_inst_req_1;
      MUX_1281_inst_ack_1<= update_ack(0);
      MUX_1281_inst: SelectSplitProtocol generic map(name => "MUX_1281_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1165_1165_delayed_1_0_1275, y => type_cast_1280_wire_constant, sel => ifx_xend_ifx_xend300_taken_1026, z => MUX_1168_1168_delayed_2_0_1282, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1289_inst
    MUX_1289_wire <= type_cast_1162_1162_delayed_1_0_1271 when (landx_xlhsx_xtrue292_ifx_xend300_taken_1229(0) /=  '0') else MUX_1168_1168_delayed_2_0_1282;
    -- flow-through select operator MUX_1290_inst
    add_outx_x2504_1291 <= type_cast_1159_1159_delayed_1_0_1267 when (ifx_xthen299_ifx_xend300_taken_1235(0) /=  '0') else MUX_1289_wire;
    MUX_1305_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1305_inst_req_0;
      MUX_1305_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1305_inst_req_1;
      MUX_1305_inst_ack_1<= update_ack(0);
      MUX_1305_inst: SelectSplitProtocol generic map(name => "MUX_1305_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1182_1182_delayed_1_0_1299, y => type_cast_1304_wire_constant, sel => ifx_xend_ifx_xend300_taken_1026, z => MUX_1185_1185_delayed_2_0_1306, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1315_inst
    MUX_1315_wire <= type_cast_1179_1179_delayed_3_0_1295 when (landx_xlhsx_xtrue292_ifx_xend300_taken_1229(0) /=  '0') else MUX_1185_1185_delayed_2_0_1306;
    -- flow-through select operator MUX_1316_inst
    count_inp1x_x2_1317 <= type_cast_1311_wire_constant when (ifx_xthen299_ifx_xend300_taken_1235(0) /=  '0') else MUX_1315_wire;
    MUX_1331_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1331_inst_req_0;
      MUX_1331_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1331_inst_req_1;
      MUX_1331_inst_ack_1<= update_ack(0);
      MUX_1331_inst: SelectSplitProtocol generic map(name => "MUX_1331_inst", data_width => 16, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1199_1199_delayed_2_0_1325, y => type_cast_1330_wire_constant, sel => ifx_xend_ifx_xend300_taken_1026, z => MUX_1202_1202_delayed_2_0_1332, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1341_inst
    MUX_1341_wire <= type_cast_1196_1196_delayed_1_0_1321 when (landx_xlhsx_xtrue292_ifx_xend300_taken_1229(0) /=  '0') else MUX_1202_1202_delayed_2_0_1332;
    -- flow-through select operator MUX_1342_inst
    count_inp2x_x2_1343 <= type_cast_1337_wire_constant when (ifx_xthen299_ifx_xend300_taken_1235(0) /=  '0') else MUX_1341_wire;
    -- flow-through select operator MUX_1522_inst
    tmp475_1523 <= xx_xop_1516 when (tmp472_1500(0) /=  '0') else type_cast_1521_wire_constant;
    -- flow-through select operator MUX_373_inst
    tmp500_374 <= xx_xop503_367 when (tmp496_351(0) /=  '0') else type_cast_372_wire_constant;
    -- flow-through select operator MUX_590_inst
    tmp487_591 <= xx_xop502_584 when (tmp483_568(0) /=  '0') else type_cast_589_wire_constant;
    -- flow-through select operator MUX_963_inst
    MUX_963_wire <= type_cast_933_933_delayed_1_0_954 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_962_wire_constant;
    -- flow-through select operator MUX_964_inst
    add_outx_x0_965 <= type_cast_958_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_963_wire;
    -- flow-through select operator MUX_978_inst
    MUX_978_wire <= type_cast_945_945_delayed_1_0_969 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_977_wire_constant;
    -- flow-through select operator MUX_979_inst
    add_inp1x_x0_980 <= type_cast_973_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_978_wire;
    -- flow-through select operator MUX_993_inst
    MUX_993_wire <= type_cast_957_957_delayed_1_0_984 when (whilex_xbody_ifx_xend_taken_860(0) /=  '0') else type_cast_992_wire_constant;
    -- flow-through select operator MUX_994_inst
    count_inp1x_x0_995 <= type_cast_988_wire when (ifx_xthen_ifx_xend_taken_945(0) /=  '0') else MUX_993_wire;
    W_add_inp1x_x1_866_delayed_1_0_864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp1x_x1_866_delayed_1_0_864_inst_req_0;
      W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp1x_x1_866_delayed_1_0_864_inst_req_1;
      W_add_inp1x_x1_866_delayed_1_0_864_inst_ack_1<= rack(0);
      W_add_inp1x_x1_866_delayed_1_0_864_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp1x_x1_866_delayed_1_0_864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp1x_x1_866_delayed_1_0_866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp1x_x1_907_delayed_1_0_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp1x_x1_907_delayed_1_0_923_inst_req_0;
      W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp1x_x1_907_delayed_1_0_923_inst_req_1;
      W_add_inp1x_x1_907_delayed_1_0_923_inst_ack_1<= rack(0);
      W_add_inp1x_x1_907_delayed_1_0_923_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp1x_x1_907_delayed_1_0_923_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp1x_x1_907_delayed_1_0_925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp2x_x1_1015_delayed_3_0_1067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_0;
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp2x_x1_1015_delayed_3_0_1067_inst_req_1;
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst_ack_1<= rack(0);
      W_add_inp2x_x1_1015_delayed_3_0_1067_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp2x_x1_1015_delayed_3_0_1067_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp2x_x1_1015_delayed_3_0_1069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_inp2x_x1_1056_delayed_3_0_1126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_0;
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_0<= wack(0);
      rreq(0) <= W_add_inp2x_x1_1056_delayed_3_0_1126_inst_req_1;
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst_ack_1<= rack(0);
      W_add_inp2x_x1_1056_delayed_3_0_1126_inst : InterlockBuffer generic map ( -- 
        name => "W_add_inp2x_x1_1056_delayed_3_0_1126_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_inp2x_x1_1056_delayed_3_0_1128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x0_1032_delayed_2_0_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x0_1032_delayed_2_0_1090_inst_req_0;
      W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x0_1032_delayed_2_0_1090_inst_req_1;
      W_add_outx_x0_1032_delayed_2_0_1090_inst_ack_1<= rack(0);
      W_add_outx_x0_1032_delayed_2_0_1090_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x0_1032_delayed_2_0_1090_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x0_1032_delayed_2_0_1092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x0_1063_delayed_2_0_1136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x0_1063_delayed_2_0_1136_inst_req_0;
      W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x0_1063_delayed_2_0_1136_inst_req_1;
      W_add_outx_x0_1063_delayed_2_0_1136_inst_ack_1<= rack(0);
      W_add_outx_x0_1063_delayed_2_0_1136_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x0_1063_delayed_2_0_1136_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x0_1063_delayed_2_0_1138,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x1_883_delayed_1_0_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x1_883_delayed_1_0_887_inst_req_0;
      W_add_outx_x1_883_delayed_1_0_887_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x1_883_delayed_1_0_887_inst_req_1;
      W_add_outx_x1_883_delayed_1_0_887_inst_ack_1<= rack(0);
      W_add_outx_x1_883_delayed_1_0_887_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x1_883_delayed_1_0_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x1_883_delayed_1_0_889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x1_914_delayed_1_0_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x1_914_delayed_1_0_933_inst_req_0;
      W_add_outx_x1_914_delayed_1_0_933_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x1_914_delayed_1_0_933_inst_req_1;
      W_add_outx_x1_914_delayed_1_0_933_inst_ack_1<= rack(0);
      W_add_outx_x1_914_delayed_1_0_933_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x1_914_delayed_1_0_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x1_914_delayed_1_0_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx252_894_delayed_6_0_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx252_894_delayed_6_0_905_inst_req_0;
      W_arrayidx252_894_delayed_6_0_905_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx252_894_delayed_6_0_905_inst_req_1;
      W_arrayidx252_894_delayed_6_0_905_inst_ack_1<= rack(0);
      W_arrayidx252_894_delayed_6_0_905_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx252_894_delayed_6_0_905_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx252_901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx252_894_delayed_6_0_907,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx278_1043_delayed_6_0_1108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx278_1043_delayed_6_0_1108_inst_req_0;
      W_arrayidx278_1043_delayed_6_0_1108_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx278_1043_delayed_6_0_1108_inst_req_1;
      W_arrayidx278_1043_delayed_6_0_1108_inst_ack_1<= rack(0);
      W_arrayidx278_1043_delayed_6_0_1108_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx278_1043_delayed_6_0_1108_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx278_1104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx278_1043_delayed_6_0_1110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp1x_x1_900_delayed_1_0_913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp1x_x1_900_delayed_1_0_913_inst_req_0;
      W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp1x_x1_900_delayed_1_0_913_inst_req_1;
      W_count_inp1x_x1_900_delayed_1_0_913_inst_ack_1<= rack(0);
      W_count_inp1x_x1_900_delayed_1_0_913_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp1x_x1_900_delayed_1_0_913_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp1x_x1_900_delayed_1_0_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp2x_x1_1049_delayed_3_0_1116_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_0;
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp2x_x1_1049_delayed_3_0_1116_inst_req_1;
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst_ack_1<= rack(0);
      W_count_inp2x_x1_1049_delayed_3_0_1116_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp2x_x1_1049_delayed_3_0_1116_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp2x_x1_1049_delayed_3_0_1118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_inp2x_x1_990_delayed_2_0_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_0;
      W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_0<= wack(0);
      rreq(0) <= W_count_inp2x_x1_990_delayed_2_0_1030_inst_req_1;
      W_count_inp2x_x1_990_delayed_2_0_1030_inst_ack_1<= rack(0);
      W_count_inp2x_x1_990_delayed_2_0_1030_inst : InterlockBuffer generic map ( -- 
        name => "W_count_inp2x_x1_990_delayed_2_0_1030_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_inp2x_x1_990_delayed_2_0_1032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xend300_whilex_xend_taken_1353_inst
    process(cmp305_1352) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp305_1352(0 downto 0);
      ifx_xend300_whilex_xend_taken_1355 <= tmp_var; -- 
    end process;
    W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_0;
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_req_1;
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_968_delayed_1_0_1001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_968_delayed_1_0_1003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_0;
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_req_1;
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_975_delayed_1_0_1010_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_975_delayed_1_0_1012,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_0;
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_req_1;
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_980_delayed_1_0_1018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_980_delayed_1_0_1020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_0;
      W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_req_1;
      W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst_ack_1<= rack(0);
      W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen271_exec_guard_1025_delayed_7_0_1082_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen271_exec_guard_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen271_exec_guard_1025_delayed_7_0_1084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_0;
      W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_req_1;
      W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst_ack_1<= rack(0);
      W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen271_exec_guard_1042_delayed_13_0_1105_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen271_exec_guard_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen271_exec_guard_1042_delayed_13_0_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen271_exec_guard_1064_inst
    process(landx_xlhsx_xtrue_ifx_xthen271_taken_1054) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue_ifx_xthen271_taken_1054(0 downto 0);
      ifx_xthen271_exec_guard_1066 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen271_landx_xlhsx_xtrue292_taken_1146_inst
    process(ifx_xthen271_exec_guard_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen271_exec_guard_1066(0 downto 0);
      ifx_xthen271_landx_xlhsx_xtrue292_taken_1148 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen299_exec_guard_1230_inst
    process(landx_xlhsx_xtrue292_ifx_xthen299_taken_1220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue292_ifx_xthen299_taken_1220(0 downto 0);
      ifx_xthen299_exec_guard_1232 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen299_ifx_xend300_taken_1233_inst
    process(ifx_xthen299_exec_guard_1232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen299_exec_guard_1232(0 downto 0);
      ifx_xthen299_ifx_xend300_taken_1235 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen_exec_guard_861_inst
    process(whilex_xbody_ifx_xthen_taken_856) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xthen_taken_856(0 downto 0);
      ifx_xthen_exec_guard_863 <= tmp_var; -- 
    end process;
    W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_0;
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_req_1;
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst_ack_1<= rack(0);
      W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_exec_guard_876_delayed_7_0_879_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_exec_guard_863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_exec_guard_876_delayed_7_0_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_0;
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_req_1;
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst_ack_1<= rack(0);
      W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_exec_guard_893_delayed_13_0_902_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_exec_guard_863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_exec_guard_893_delayed_13_0_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen_ifx_xend_taken_943_inst
    process(ifx_xthen_exec_guard_863) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen_exec_guard_863(0 downto 0);
      ifx_xthen_ifx_xend_taken_945 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_0;
      W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_req_1;
      W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue292_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue292_exec_guard_1117_delayed_1_0_1206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_0;
      W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_req_1;
      W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1213_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue292_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_0;
      W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_req_1;
      W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1221_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue292_exec_guard_1153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1047_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1055_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_landx_xlhsx_xtrue_exec_guard_1027_inst
    process(ifx_xend_landx_xlhsx_xtrue_taken_1017) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend_landx_xlhsx_xtrue_taken_1017(0 downto 0);
      landx_xlhsx_xtrue_exec_guard_1029 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_0;
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_req_1;
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue_exec_guard_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue_exec_guard_993_delayed_1_0_1040,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_ifx_xthen_taken_854_inst
    process(cmp244_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp244_853(0 downto 0);
      whilex_xbody_ifx_xthen_taken_856 <= tmp_var; -- 
    end process;
    addr_of_1080_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1080_final_reg_req_0;
      addr_of_1080_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1080_final_reg_req_1;
      addr_of_1080_final_reg_ack_1<= rack(0);
      addr_of_1080_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1080_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1079_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx274_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1103_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1103_final_reg_req_0;
      addr_of_1103_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1103_final_reg_req_1;
      addr_of_1103_final_reg_ack_1<= rack(0);
      addr_of_1103_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1103_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1102_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx278_1104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1539_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1539_final_reg_req_0;
      addr_of_1539_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1539_final_reg_req_1;
      addr_of_1539_final_reg_ack_1<= rack(0);
      addr_of_1539_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1539_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1538_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx388_1540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_390_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_390_final_reg_req_0;
      addr_of_390_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_390_final_reg_req_1;
      addr_of_390_final_reg_ack_1<= rack(0);
      addr_of_390_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_390_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_389_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_607_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_607_final_reg_req_0;
      addr_of_607_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_607_final_reg_req_1;
      addr_of_607_final_reg_ack_1<= rack(0);
      addr_of_607_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_607_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_606_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx227_608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_877_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_877_final_reg_req_0;
      addr_of_877_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_877_final_reg_req_1;
      addr_of_877_final_reg_ack_1<= rack(0);
      addr_of_877_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_877_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_876_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx248_878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_900_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_900_final_reg_req_0;
      addr_of_900_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_900_final_reg_req_1;
      addr_of_900_final_reg_ack_1<= rack(0);
      addr_of_900_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_900_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_899_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx252_901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1036_inst_req_0;
      type_cast_1036_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1036_inst_req_1;
      type_cast_1036_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue_exec_guard_1029(0);
      type_cast_1036_inst_gI: SplitGuardInterface generic map(name => "type_cast_1036_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1036_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_990_delayed_2_0_1032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv266_1037,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_105_inst_req_0;
      type_cast_105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_105_inst_req_1;
      type_cast_105_inst_ack_1<= rack(0);
      type_cast_105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_102,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1073_inst_req_0;
      type_cast_1073_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1073_inst_req_1;
      type_cast_1073_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen271_exec_guard_1066(0);
      type_cast_1073_inst_gI: SplitGuardInterface generic map(name => "type_cast_1073_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1073_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_1015_delayed_3_0_1069,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom273_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1096_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1096_inst_req_0;
      type_cast_1096_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1096_inst_req_1;
      type_cast_1096_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen271_exec_guard_1066(0);
      type_cast_1096_inst_gI: SplitGuardInterface generic map(name => "type_cast_1096_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1096_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1096_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_1032_delayed_2_0_1092,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom277_1097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1156_inst_req_0;
      type_cast_1156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1156_inst_req_1;
      type_cast_1156_inst_ack_1<= rack(0);
      type_cast_1156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1156_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1082_1082_delayed_2_0_1157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1161_inst
    process(inc284_1145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc284_1145(15 downto 0);
      type_cast_1161_wire <= tmp_var; -- 
    end process;
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1094_1094_delayed_3_0_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1176_inst
    process(inc282_1135) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc282_1135(15 downto 0);
      type_cast_1176_wire <= tmp_var; -- 
    end process;
    type_cast_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1186_inst_req_0;
      type_cast_1186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1186_inst_req_1;
      type_cast_1186_inst_ack_1<= rack(0);
      type_cast_1186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1186_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1106_1106_delayed_3_0_1187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_118_inst_req_0;
      type_cast_118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_118_inst_req_1;
      type_cast_118_inst_ack_1<= rack(0);
      type_cast_118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1191_inst
    process(inc280_1125) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc280_1125(15 downto 0);
      type_cast_1191_wire <= tmp_var; -- 
    end process;
    type_cast_1202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1202_inst_req_0;
      type_cast_1202_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1202_inst_req_1;
      type_cast_1202_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue292_exec_guard_1153(0);
      type_cast_1202_inst_gI: SplitGuardInterface generic map(name => "type_cast_1202_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1202_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x0x_xph_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv294_1203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0x_xph_1183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1143_1143_delayed_1_0_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1242_inst_req_0;
      type_cast_1242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1242_inst_req_1;
      type_cast_1242_inst_ack_1<= rack(0);
      type_cast_1242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1242_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0x_xph_1183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1146_1146_delayed_1_0_1243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1246_inst_req_0;
      type_cast_1246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1246_inst_req_1;
      type_cast_1246_inst_ack_1<= rack(0);
      type_cast_1246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1246_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x1_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1149_1149_delayed_2_0_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2x_xph_1168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1159_1159_delayed_1_0_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1270_inst_req_0;
      type_cast_1270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1270_inst_req_1;
      type_cast_1270_inst_ack_1<= rack(0);
      type_cast_1270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1270_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2x_xph_1168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1162_1162_delayed_1_0_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1274_inst_req_0;
      type_cast_1274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1274_inst_req_1;
      type_cast_1274_inst_ack_1<= rack(0);
      type_cast_1274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1165_1165_delayed_1_0_1275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1294_inst_req_0;
      type_cast_1294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1294_inst_req_1;
      type_cast_1294_inst_ack_1<= rack(0);
      type_cast_1294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1294_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1179_1179_delayed_3_0_1295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1298_inst_req_0;
      type_cast_1298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1298_inst_req_1;
      type_cast_1298_inst_ack_1<= rack(0);
      type_cast_1298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1182_1182_delayed_1_0_1299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_130_inst_req_0;
      type_cast_130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_130_inst_req_1;
      type_cast_130_inst_ack_1<= rack(0);
      type_cast_130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x0x_xph_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1196_1196_delayed_1_0_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1324_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1324_inst_req_0;
      type_cast_1324_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1324_inst_req_1;
      type_cast_1324_inst_ack_1<= rack(0);
      type_cast_1324_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1324_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x1_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1199_1199_delayed_2_0_1325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2504_1291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv302_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1367_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv234_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1375_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1385_inst_req_0;
      type_cast_1385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1385_inst_req_1;
      type_cast_1385_inst_ack_1<= rack(0);
      type_cast_1385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1395_inst_req_0;
      type_cast_1395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1395_inst_req_1;
      type_cast_1395_inst_ack_1<= rack(0);
      type_cast_1395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_1392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_1396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1405_inst_req_0;
      type_cast_1405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1405_inst_req_1;
      type_cast_1405_inst_ack_1<= rack(0);
      type_cast_1405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_1402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_1406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1415_inst_req_0;
      type_cast_1415_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1415_inst_req_1;
      type_cast_1415_inst_ack_1<= rack(0);
      type_cast_1415_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1415_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_1412,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_1416,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1435_inst_req_0;
      type_cast_1435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1435_inst_req_1;
      type_cast_1435_inst_ack_1<= rack(0);
      type_cast_1435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_143_inst_req_0;
      type_cast_143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_143_inst_req_1;
      type_cast_143_inst_ack_1<= rack(0);
      type_cast_143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1445_inst_req_0;
      type_cast_1445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1445_inst_req_1;
      type_cast_1445_inst_ack_1<= rack(0);
      type_cast_1445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr350_1442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv353_1446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1455_inst_req_0;
      type_cast_1455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1455_inst_req_1;
      type_cast_1455_inst_ack_1<= rack(0);
      type_cast_1455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr356_1452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv359_1456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1509_inst_req_0;
      type_cast_1509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1509_inst_req_1;
      type_cast_1509_inst_ack_1<= rack(0);
      type_cast_1509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp471x_xop_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_79_1510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1532_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1532_inst_req_0;
      type_cast_1532_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1532_inst_req_1;
      type_cast_1532_inst_ack_1<= rack(0);
      type_cast_1532_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1532_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1532_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1547_inst_req_0;
      type_cast_1547_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1547_inst_req_1;
      type_cast_1547_inst_ack_1<= rack(0);
      type_cast_1547_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1547_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_1544,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv393_1548,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1557_inst_req_0;
      type_cast_1557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1557_inst_req_1;
      type_cast_1557_inst_ack_1<= rack(0);
      type_cast_1557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr396_1554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_1558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_156,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1567_inst_req_0;
      type_cast_1567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1567_inst_req_1;
      type_cast_1567_inst_ack_1<= rack(0);
      type_cast_1567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr402_1564,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv405_1568,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1577_inst_req_0;
      type_cast_1577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1577_inst_req_1;
      type_cast_1577_inst_ack_1<= rack(0);
      type_cast_1577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr408_1574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1587_inst_req_0;
      type_cast_1587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1587_inst_req_1;
      type_cast_1587_inst_ack_1<= rack(0);
      type_cast_1587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1597_inst_req_0;
      type_cast_1597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1597_inst_req_1;
      type_cast_1597_inst_ack_1<= rack(0);
      type_cast_1597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr420_1594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv423_1598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1607_inst_req_0;
      type_cast_1607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1607_inst_req_1;
      type_cast_1607_inst_ack_1<= rack(0);
      type_cast_1607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr426_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv429_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1617_inst_req_0;
      type_cast_1617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1617_inst_req_1;
      type_cast_1617_inst_ack_1<= rack(0);
      type_cast_1617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr432_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv435_1618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_168_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_168_inst_req_0;
      type_cast_168_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_168_inst_req_1;
      type_cast_168_inst_ack_1<= rack(0);
      type_cast_168_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_168_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_169,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_180_inst_req_0;
      type_cast_180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_180_inst_req_1;
      type_cast_180_inst_ack_1<= rack(0);
      type_cast_180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_193_inst_req_0;
      type_cast_193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_193_inst_req_1;
      type_cast_193_inst_ack_1<= rack(0);
      type_cast_193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_230_inst_req_0;
      type_cast_230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_230_inst_req_1;
      type_cast_230_inst_ack_1<= rack(0);
      type_cast_230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_243_inst_req_0;
      type_cast_243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_243_inst_req_1;
      type_cast_243_inst_ack_1<= rack(0);
      type_cast_243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_30_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_30_inst_req_0;
      type_cast_30_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_30_inst_req_1;
      type_cast_30_inst_ack_1<= rack(0);
      type_cast_30_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_30_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_26,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_31,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_360_inst_req_0;
      type_cast_360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_360_inst_req_1;
      type_cast_360_inst_ack_1<= rack(0);
      type_cast_360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp495x_xop_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_383_inst_req_0;
      type_cast_383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_383_inst_req_1;
      type_cast_383_inst_ack_1<= rack(0);
      type_cast_383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext490_534,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_383_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_397_inst_req_0;
      type_cast_397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_397_inst_req_1;
      type_cast_397_inst_ack_1<= rack(0);
      type_cast_397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_410_inst_req_0;
      type_cast_410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_410_inst_req_1;
      type_cast_410_inst_ack_1<= rack(0);
      type_cast_410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_407,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_428_inst_req_0;
      type_cast_428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_428_inst_req_1;
      type_cast_428_inst_ack_1<= rack(0);
      type_cast_428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_43_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_43_inst_req_0;
      type_cast_43_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_43_inst_req_1;
      type_cast_43_inst_ack_1<= rack(0);
      type_cast_43_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_43_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_40,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_44,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_446_inst_req_0;
      type_cast_446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_446_inst_req_1;
      type_cast_446_inst_ack_1<= rack(0);
      type_cast_446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call140_443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_464_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_464_inst_req_0;
      type_cast_464_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_464_inst_req_1;
      type_cast_464_inst_ack_1<= rack(0);
      type_cast_464_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_464_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call146_461,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_482_inst_req_0;
      type_cast_482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_482_inst_req_1;
      type_cast_482_inst_ack_1<= rack(0);
      type_cast_482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_500_inst_req_0;
      type_cast_500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_500_inst_req_1;
      type_cast_500_inst_ack_1<= rack(0);
      type_cast_500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call158_497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_518_inst_req_0;
      type_cast_518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_518_inst_req_1;
      type_cast_518_inst_ack_1<= rack(0);
      type_cast_518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_55_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_55_inst_req_0;
      type_cast_55_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_55_inst_req_1;
      type_cast_55_inst_ack_1<= rack(0);
      type_cast_55_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_55_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_52,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_56,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp482x_xop_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_32_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_600_inst_req_0;
      type_cast_600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_600_inst_req_1;
      type_cast_600_inst_ack_1<= rack(0);
      type_cast_600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_600_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_614_inst_req_1;
      type_cast_614_inst_ack_1<= rack(0);
      type_cast_614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_627_inst_req_0;
      type_cast_627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_627_inst_req_1;
      type_cast_627_inst_ack_1<= rack(0);
      type_cast_627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call184_624,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_628,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_645_inst_req_0;
      type_cast_645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_645_inst_req_1;
      type_cast_645_inst_ack_1<= rack(0);
      type_cast_645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call190_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_663_inst_req_0;
      type_cast_663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_663_inst_req_1;
      type_cast_663_inst_ack_1<= rack(0);
      type_cast_663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call196_660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_681_inst_req_0;
      type_cast_681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_681_inst_req_1;
      type_cast_681_inst_ack_1<= rack(0);
      type_cast_681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call202_678,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv204_682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_68_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_68_inst_req_0;
      type_cast_68_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_68_inst_req_1;
      type_cast_68_inst_ack_1<= rack(0);
      type_cast_68_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_68_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_65,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_69,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call208_696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_717_inst_req_0;
      type_cast_717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_717_inst_req_1;
      type_cast_717_inst_ack_1<= rack(0);
      type_cast_717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call214_714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_735_inst_req_0;
      type_cast_735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_735_inst_req_1;
      type_cast_735_inst_ack_1<= rack(0);
      type_cast_735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call220_732,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv222_736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_80_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_80_inst_req_0;
      type_cast_80_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_80_inst_req_1;
      type_cast_80_inst_ack_1<= rack(0);
      type_cast_80_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_80_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_77,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_81,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x2504_1291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_822_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_827_inst_req_0;
      type_cast_827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_827_inst_req_1;
      type_cast_827_inst_ack_1<= rack(0);
      type_cast_827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_827_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x0_980,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_827_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp2x_x0506_1263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_837_inst_req_0;
      type_cast_837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_837_inst_req_1;
      type_cast_837_inst_ack_1<= rack(0);
      type_cast_837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_837_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x2_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_837_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp2x_x2_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_842_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_870_inst_req_0;
      type_cast_870_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_870_inst_req_1;
      type_cast_870_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen_exec_guard_863(0);
      type_cast_870_inst_gI: SplitGuardInterface generic map(name => "type_cast_870_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_866_delayed_1_0_866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom247_871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_893_inst_req_0;
      type_cast_893_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_893_inst_req_1;
      type_cast_893_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen_exec_guard_863(0);
      type_cast_893_inst_gI: SplitGuardInterface generic map(name => "type_cast_893_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_883_delayed_1_0_889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom251_894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_93_inst_req_0;
      type_cast_93_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_93_inst_req_1;
      type_cast_93_inst_ack_1<= rack(0);
      type_cast_93_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_93_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_90,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_94,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_953_inst_req_0;
      type_cast_953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_953_inst_req_1;
      type_cast_953_inst_ack_1<= rack(0);
      type_cast_953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_933_933_delayed_1_0_954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_958_inst
    process(inc258_942) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc258_942(15 downto 0);
      type_cast_958_wire <= tmp_var; -- 
    end process;
    type_cast_968_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_968_inst_req_0;
      type_cast_968_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_968_inst_req_1;
      type_cast_968_inst_ack_1<= rack(0);
      type_cast_968_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_968_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_inp1x_x1_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_945_945_delayed_1_0_969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_973_inst
    process(inc256_932) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc256_932(15 downto 0);
      type_cast_973_wire <= tmp_var; -- 
    end process;
    type_cast_983_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_983_inst_req_0;
      type_cast_983_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_983_inst_req_1;
      type_cast_983_inst_ack_1<= rack(0);
      type_cast_983_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_983_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x1_834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_957_957_delayed_1_0_984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_988_inst
    process(inc254_922) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := inc254_922(15 downto 0);
      type_cast_988_wire <= tmp_var; -- 
    end process;
    type_cast_999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_999_inst_req_0;
      type_cast_999_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_999_inst_req_1;
      type_cast_999_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend_exec_guard_950(0);
      type_cast_999_inst_gI: SplitGuardInterface generic map(name => "type_cast_999_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_999_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_inp1x_x0_995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv260_1000,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1079_index_1_rename
    process(R_idxprom273_1078_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom273_1078_resized;
      ov(13 downto 0) := iv;
      R_idxprom273_1078_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_index_1_resize
    process(idxprom273_1074) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom273_1074;
      ov := iv(13 downto 0);
      R_idxprom273_1078_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_root_address_inst
    process(array_obj_ref_1079_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1079_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_index_1_rename
    process(R_idxprom277_1101_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom277_1101_resized;
      ov(13 downto 0) := iv;
      R_idxprom277_1101_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_index_1_resize
    process(idxprom277_1097) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom277_1097;
      ov := iv(13 downto 0);
      R_idxprom277_1101_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1102_root_address_inst
    process(array_obj_ref_1102_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1102_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1102_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_index_1_rename
    process(R_indvar_1537_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1537_resized;
      ov(13 downto 0) := iv;
      R_indvar_1537_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_index_1_resize
    process(indvar_1526) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1526;
      ov := iv(13 downto 0);
      R_indvar_1537_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1538_root_address_inst
    process(array_obj_ref_1538_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1538_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1538_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_389_index_1_rename
    process(R_indvar489_388_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar489_388_resized;
      ov(13 downto 0) := iv;
      R_indvar489_388_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_389_index_1_resize
    process(indvar489_377) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar489_377;
      ov := iv(13 downto 0);
      R_indvar489_388_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_389_root_address_inst
    process(array_obj_ref_389_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_389_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_389_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_606_index_1_rename
    process(R_indvar476_605_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_605_resized;
      ov(13 downto 0) := iv;
      R_indvar476_605_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_606_index_1_resize
    process(indvar476_594) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_594;
      ov := iv(13 downto 0);
      R_indvar476_605_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_606_root_address_inst
    process(array_obj_ref_606_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_606_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_606_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_rename
    process(R_idxprom247_875_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom247_875_resized;
      ov(13 downto 0) := iv;
      R_idxprom247_875_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_resize
    process(idxprom247_871) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom247_871;
      ov := iv(13 downto 0);
      R_idxprom247_875_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_root_address_inst
    process(array_obj_ref_876_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_876_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_876_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_index_1_rename
    process(R_idxprom251_898_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom251_898_resized;
      ov(13 downto 0) := iv;
      R_idxprom251_898_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_index_1_resize
    process(idxprom251_894) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom251_894;
      ov := iv(13 downto 0);
      R_idxprom251_898_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_899_root_address_inst
    process(array_obj_ref_899_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_899_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_899_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_addr_0
    process(ptr_deref_1088_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_base_resize
    process(arrayidx274_1081) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx274_1081;
      ov := iv(13 downto 0);
      ptr_deref_1088_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_gather_scatter
    process(ptr_deref_1088_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_data_0;
      ov(63 downto 0) := iv;
      tmp275_1089 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1088_root_address_inst
    process(ptr_deref_1088_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1088_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1088_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_addr_0
    process(ptr_deref_1113_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1113_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_base_resize
    process(arrayidx278_1043_delayed_6_0_1110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx278_1043_delayed_6_0_1110;
      ov := iv(13 downto 0);
      ptr_deref_1113_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_gather_scatter
    process(tmp275_1089) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp275_1089;
      ov(63 downto 0) := iv;
      ptr_deref_1113_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_root_address_inst
    process(ptr_deref_1113_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1113_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_addr_0
    process(ptr_deref_1543_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1543_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_base_resize
    process(arrayidx388_1540) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx388_1540;
      ov := iv(13 downto 0);
      ptr_deref_1543_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_gather_scatter
    process(ptr_deref_1543_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_data_0;
      ov(63 downto 0) := iv;
      tmp389_1544 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1543_root_address_inst
    process(ptr_deref_1543_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1543_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1543_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_addr_0
    process(ptr_deref_526_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_526_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_526_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_base_resize
    process(arrayidx_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_391;
      ov := iv(13 downto 0);
      ptr_deref_526_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_gather_scatter
    process(add167_524) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add167_524;
      ov(63 downto 0) := iv;
      ptr_deref_526_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_526_root_address_inst
    process(ptr_deref_526_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_526_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_526_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_addr_0
    process(ptr_deref_743_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_743_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_743_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_base_resize
    process(arrayidx227_608) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx227_608;
      ov := iv(13 downto 0);
      ptr_deref_743_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_gather_scatter
    process(add223_741) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add223_741;
      ov(63 downto 0) := iv;
      ptr_deref_743_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_743_root_address_inst
    process(ptr_deref_743_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_743_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_743_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_addr_0
    process(ptr_deref_885_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_885_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_base_resize
    process(arrayidx248_878) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx248_878;
      ov := iv(13 downto 0);
      ptr_deref_885_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_gather_scatter
    process(ptr_deref_885_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_data_0;
      ov(63 downto 0) := iv;
      tmp249_886 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_885_root_address_inst
    process(ptr_deref_885_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_885_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_885_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_addr_0
    process(ptr_deref_910_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_910_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_910_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_base_resize
    process(arrayidx252_894_delayed_6_0_907) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx252_894_delayed_6_0_907;
      ov := iv(13 downto 0);
      ptr_deref_910_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_gather_scatter
    process(tmp249_886) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp249_886;
      ov(63 downto 0) := iv;
      ptr_deref_910_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_910_root_address_inst
    process(ptr_deref_910_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_910_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_910_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_817_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1358_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_817_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_817_branch_req_0,
          ack0 => do_while_stmt_817_branch_ack_0,
          ack1 => do_while_stmt_817_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1359_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend300_whilex_xend_taken_1355;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1359_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1359_branch_req_0,
          ack0 => if_stmt_1359_branch_ack_0,
          ack1 => if_stmt_1359_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1488_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp381460_1487;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1488_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1488_branch_req_0,
          ack0 => if_stmt_1488_branch_ack_0,
          ack1 => if_stmt_1488_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1654_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1653;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1654_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1654_branch_req_0,
          ack0 => if_stmt_1654_branch_ack_0,
          ack1 => if_stmt_1654_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_308_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp467_307;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_308_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_308_branch_req_0,
          ack0 => if_stmt_308_branch_ack_0,
          ack1 => if_stmt_308_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_323_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp175463_322;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_323_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_323_branch_req_0,
          ack0 => if_stmt_323_branch_ack_0,
          ack1 => if_stmt_323_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_540_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_539;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_540_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_540_branch_req_0,
          ack0 => if_stmt_540_branch_ack_0,
          ack1 => if_stmt_540_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_757_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_756;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_757_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_757_branch_req_0,
          ack0 => if_stmt_757_branch_ack_0,
          ack1 => if_stmt_757_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1124_inst
    process(count_inp2x_x1_1049_delayed_3_0_1118) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp2x_x1_1049_delayed_3_0_1118, type_cast_1123_wire_constant, tmp_var);
      inc280_1125 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1134_inst
    process(add_inp2x_x1_1056_delayed_3_0_1128) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp2x_x1_1056_delayed_3_0_1128, type_cast_1133_wire_constant, tmp_var);
      inc282_1135 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1144_inst
    process(add_outx_x0_1063_delayed_2_0_1138) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_outx_x0_1063_delayed_2_0_1138, type_cast_1143_wire_constant, tmp_var);
      inc284_1145 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_921_inst
    process(count_inp1x_x1_900_delayed_1_0_915) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp1x_x1_900_delayed_1_0_915, type_cast_920_wire_constant, tmp_var);
      inc254_922 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_931_inst
    process(add_inp1x_x1_907_delayed_1_0_925) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp1x_x1_907_delayed_1_0_925, type_cast_930_wire_constant, tmp_var);
      inc256_932 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_941_inst
    process(add_outx_x1_914_delayed_1_0_935) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_outx_x1_914_delayed_1_0_935, type_cast_940_wire_constant, tmp_var);
      inc258_942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1505_inst
    process(shr304_787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr304_787, type_cast_1504_wire_constant, tmp_var);
      tmp471x_xop_1506 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_356_inst
    process(tmp495_345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp495_345, type_cast_355_wire_constant, tmp_var);
      tmp495x_xop_357 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_573_inst
    process(tmp482_562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp482_562, type_cast_572_wire_constant, tmp_var);
      tmp482x_xop_574 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1515_inst
    process(iNsTr_79_1510) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_79_1510, type_cast_1514_wire_constant, tmp_var);
      xx_xop_1516 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1647_inst
    process(indvar_1526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1526, type_cast_1646_wire_constant, tmp_var);
      indvarx_xnext_1648 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_366_inst
    process(iNsTr_19_361) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_19_361, type_cast_365_wire_constant, tmp_var);
      xx_xop503_367 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_533_inst
    process(indvar489_377) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar489_377, type_cast_532_wire_constant, tmp_var);
      indvarx_xnext490_534 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_583_inst
    process(iNsTr_32_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_32_578, type_cast_582_wire_constant, tmp_var);
      xx_xop502_584 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_750_inst
    process(indvar476_594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_594, type_cast_749_wire_constant, tmp_var);
      indvarx_xnext477_751 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1016_inst
    process(ifx_xend_exec_guard_975_delayed_1_0_1012, cmp263_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_975_delayed_1_0_1012, cmp263_1009, tmp_var);
      ifx_xend_landx_xlhsx_xtrue_taken_1017 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1025_inst
    process(ifx_xend_exec_guard_980_delayed_1_0_1020, NOT_u1_u1_1024_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_980_delayed_1_0_1020, NOT_u1_u1_1024_wire, tmp_var);
      ifx_xend_ifx_xend300_taken_1026 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1053_inst
    process(landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049, cmp269_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue_exec_guard_1000_delayed_1_0_1049, cmp269_1046, tmp_var);
      landx_xlhsx_xtrue_ifx_xthen271_taken_1054 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1062_inst
    process(landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057, NOT_u1_u1_1061_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue_exec_guard_1005_delayed_1_0_1057, NOT_u1_u1_1061_wire, tmp_var);
      landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1219_inst
    process(landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1215, cmp297_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue292_exec_guard_1124_delayed_1_0_1215, cmp297_1212, tmp_var);
      landx_xlhsx_xtrue292_ifx_xthen299_taken_1220 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1228_inst
    process(landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1223, NOT_u1_u1_1227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue292_exec_guard_1129_delayed_1_0_1223, NOT_u1_u1_1227_wire, tmp_var);
      landx_xlhsx_xtrue292_ifx_xend300_taken_1229 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_774_inst
    process(shr457_290) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr457_290, type_cast_773_wire_constant, tmp_var);
      conv243_775 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_780_inst
    process(shr117458_301) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr117458_301, type_cast_779_wire_constant, tmp_var);
      conv268_781 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1008_inst
    process(conv260_1000, conv243_775) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv260_1000, conv243_775, tmp_var);
      cmp263_1009 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1211_inst
    process(conv294_1203, conv268_781) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv294_1203, conv268_781, tmp_var);
      cmp297_1212 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1351_inst
    process(conv302_1347, shr304_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv302_1347, shr304_787, tmp_var);
      cmp305_1352 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1652_inst
    process(indvarx_xnext_1648, tmp475_1523) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1648, tmp475_1523, tmp_var);
      exitcond1_1653 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_538_inst
    process(indvarx_xnext490_534, tmp500_374) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext490_534, tmp500_374, tmp_var);
      exitcond2_539 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_755_inst
    process(indvarx_xnext477_751, tmp487_591) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_751, tmp487_591, tmp_var);
      exitcond_756 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_289_inst
    process(mul109_284) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul109_284, type_cast_288_wire_constant, tmp_var);
      shr457_290 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_300_inst
    process(mul116_295) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul116_295, type_cast_299_wire_constant, tmp_var);
      shr117458_301 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_344_inst
    process(tmp494_339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp494_339, type_cast_343_wire_constant, tmp_var);
      tmp495_345 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_561_inst
    process(tmp481_556) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp481_556, type_cast_560_wire_constant, tmp_var);
      tmp482_562 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_786_inst
    process(mul103_279) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul103_279, type_cast_785_wire_constant, tmp_var);
      shr304_787 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1391_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1390_wire_constant, tmp_var);
      shr320_1392 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1401_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1400_wire_constant, tmp_var);
      shr326_1402 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1411_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1410_wire_constant, tmp_var);
      shr332_1412 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1421_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1420_wire_constant, tmp_var);
      shr338_1422 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1431_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1430_wire_constant, tmp_var);
      shr344_1432 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1441_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1440_wire_constant, tmp_var);
      shr350_1442 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1451_inst
    process(sub_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1382, type_cast_1450_wire_constant, tmp_var);
      shr356_1452 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1553_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1552_wire_constant, tmp_var);
      shr396_1554 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1563_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1562_wire_constant, tmp_var);
      shr402_1564 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1573_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1572_wire_constant, tmp_var);
      shr408_1574 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1583_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1582_wire_constant, tmp_var);
      shr414_1584 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1593_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1592_wire_constant, tmp_var);
      shr420_1594 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1603_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1602_wire_constant, tmp_var);
      shr426_1604 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1613_inst
    process(tmp389_1544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp389_1544, type_cast_1612_wire_constant, tmp_var);
      shr432_1614 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_253_inst
    process(add12_74, add_49) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_74, add_49, tmp_var);
      mul_254 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_258_inst
    process(mul_254, add21_99) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_254, add21_99, tmp_var);
      mul85_259 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_263_inst
    process(add39_149, add30_124) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add39_149, add30_124, tmp_var);
      mul91_264 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_268_inst
    process(mul91_264, add48_174) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul91_264, add48_174, tmp_var);
      mul94_269 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_273_inst
    process(add66_224, add57_199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add66_224, add57_199, tmp_var);
      mul100_274 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(mul100_274, add75_249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul100_274, add75_249, tmp_var);
      mul103_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(add21_99, add12_74) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add21_99, add12_74, tmp_var);
      mul109_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_294_inst
    process(add48_174, add39_149) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add48_174, add39_149, tmp_var);
      mul116_295 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_333_inst
    process(add_49, add12_74) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_49, add12_74, tmp_var);
      tmp492_334 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_338_inst
    process(tmp492_334, add21_99) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp492_334, add21_99, tmp_var);
      tmp494_339 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_550_inst
    process(add30_124, add39_149) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add30_124, add39_149, tmp_var);
      tmp479_551 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_555_inst
    process(tmp479_551, add48_174) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp479_551, add48_174, tmp_var);
      tmp481_556 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1024_inst
    process(cmp263_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp263_1009, tmp_var);
      NOT_u1_u1_1024_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1061_inst
    process(cmp269_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp269_1046, tmp_var);
      NOT_u1_u1_1061_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1227_inst
    process(cmp297_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp297_1212, tmp_var);
      NOT_u1_u1_1227_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1358_inst
    process(cmp305_1352) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp305_1352, tmp_var);
      NOT_u1_u1_1358_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_859_inst
    process(cmp244_853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp244_853, tmp_var);
      whilex_xbody_ifx_xend_taken_860 <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1152_inst
    process(ifx_xthen271_landx_xlhsx_xtrue292_taken_1148, landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen271_landx_xlhsx_xtrue292_taken_1148, landx_xlhsx_xtrue_landx_xlhsx_xtrue292_taken_1063, tmp_var);
      landx_xlhsx_xtrue292_exec_guard_1153 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_949_inst
    process(ifx_xthen_ifx_xend_taken_945, whilex_xbody_ifx_xend_taken_860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen_ifx_xend_taken_945, whilex_xbody_ifx_xend_taken_860, tmp_var);
      ifx_xend_exec_guard_950 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_123_inst
    process(shl27_112, conv29_119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_112, conv29_119, tmp_var);
      add30_124 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_148_inst
    process(shl36_137, conv38_144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_137, conv38_144, tmp_var);
      add39_149 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_173_inst
    process(shl45_162, conv47_169) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_162, conv47_169, tmp_var);
      add48_174 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_198_inst
    process(shl54_187, conv56_194) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_187, conv56_194, tmp_var);
      add57_199 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_223_inst
    process(shl63_212, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl63_212, conv65_219, tmp_var);
      add66_224 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_248_inst
    process(shl72_237, conv74_244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl72_237, conv74_244, tmp_var);
      add75_249 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_48_inst
    process(shl_37, conv3_44) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_37, conv3_44, tmp_var);
      add_49 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_73_inst
    process(shl9_62, conv11_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_62, conv11_69, tmp_var);
      add12_74 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_98_inst
    process(shl18_87, conv20_94) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_87, conv20_94, tmp_var);
      add21_99 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_415_inst
    process(shl127_404, conv130_411) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl127_404, conv130_411, tmp_var);
      add131_416 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_433_inst
    process(shl133_422, conv136_429) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl133_422, conv136_429, tmp_var);
      add137_434 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_451_inst
    process(shl139_440, conv142_447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl139_440, conv142_447, tmp_var);
      add143_452 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_469_inst
    process(shl145_458, conv148_465) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl145_458, conv148_465, tmp_var);
      add149_470 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_487_inst
    process(shl151_476, conv154_483) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl151_476, conv154_483, tmp_var);
      add155_488 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_505_inst
    process(shl157_494, conv160_501) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl157_494, conv160_501, tmp_var);
      add161_506 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_523_inst
    process(shl163_512, conv166_519) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_512, conv166_519, tmp_var);
      add167_524 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_632_inst
    process(shl183_621, conv186_628) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl183_621, conv186_628, tmp_var);
      add187_633 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_650_inst
    process(shl189_639, conv192_646) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl189_639, conv192_646, tmp_var);
      add193_651 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_668_inst
    process(shl195_657, conv198_664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl195_657, conv198_664, tmp_var);
      add199_669 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_686_inst
    process(shl201_675, conv204_682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl201_675, conv204_682, tmp_var);
      add205_687 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_704_inst
    process(shl207_693, conv210_700) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl207_693, conv210_700, tmp_var);
      add211_705 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_722_inst
    process(shl213_711, conv216_718) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl213_711, conv216_718, tmp_var);
      add217_723 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_740_inst
    process(shl219_729, conv222_736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl219_729, conv222_736, tmp_var);
      add223_741 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_111_inst
    process(conv26_106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_106, type_cast_110_wire_constant, tmp_var);
      shl27_112 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_136_inst
    process(conv35_131) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_131, type_cast_135_wire_constant, tmp_var);
      shl36_137 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_161_inst
    process(conv44_156) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_156, type_cast_160_wire_constant, tmp_var);
      shl45_162 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_186_inst
    process(conv53_181) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_181, type_cast_185_wire_constant, tmp_var);
      shl54_187 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_211_inst
    process(conv62_206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv62_206, type_cast_210_wire_constant, tmp_var);
      shl63_212 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_236_inst
    process(conv71_231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71_231, type_cast_235_wire_constant, tmp_var);
      shl72_237 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_36_inst
    process(conv1_31) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_31, type_cast_35_wire_constant, tmp_var);
      shl_37 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_61_inst
    process(conv8_56) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_56, type_cast_60_wire_constant, tmp_var);
      shl9_62 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_86_inst
    process(conv17_81) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_81, type_cast_85_wire_constant, tmp_var);
      shl18_87 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_403_inst
    process(conv125_398) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv125_398, type_cast_402_wire_constant, tmp_var);
      shl127_404 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_421_inst
    process(add131_416) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add131_416, type_cast_420_wire_constant, tmp_var);
      shl133_422 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_439_inst
    process(add137_434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add137_434, type_cast_438_wire_constant, tmp_var);
      shl139_440 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_457_inst
    process(add143_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add143_452, type_cast_456_wire_constant, tmp_var);
      shl145_458 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_475_inst
    process(add149_470) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add149_470, type_cast_474_wire_constant, tmp_var);
      shl151_476 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_493_inst
    process(add155_488) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add155_488, type_cast_492_wire_constant, tmp_var);
      shl157_494 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_511_inst
    process(add161_506) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add161_506, type_cast_510_wire_constant, tmp_var);
      shl163_512 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_620_inst
    process(conv181_615) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv181_615, type_cast_619_wire_constant, tmp_var);
      shl183_621 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_638_inst
    process(add187_633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add187_633, type_cast_637_wire_constant, tmp_var);
      shl189_639 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_656_inst
    process(add193_651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add193_651, type_cast_655_wire_constant, tmp_var);
      shl195_657 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_674_inst
    process(add199_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add199_669, type_cast_673_wire_constant, tmp_var);
      shl201_675 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_692_inst
    process(add205_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add205_687, type_cast_691_wire_constant, tmp_var);
      shl207_693 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_710_inst
    process(add211_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add211_705, type_cast_709_wire_constant, tmp_var);
      shl213_711 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_728_inst
    process(add217_723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add217_723, type_cast_727_wire_constant, tmp_var);
      shl219_729 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1381_inst
    process(conv311_1377, conv234_1369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv311_1377, conv234_1369, tmp_var);
      sub_1382 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1486_inst
    process(mul103_279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul103_279, type_cast_1485_wire_constant, tmp_var);
      cmp381460_1487 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1499_inst
    process(shr304_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr304_787, type_cast_1498_wire_constant, tmp_var);
      tmp472_1500 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_306_inst
    process(mul85_259) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul85_259, type_cast_305_wire_constant, tmp_var);
      cmp467_307 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_321_inst
    process(mul94_269) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul94_269, type_cast_320_wire_constant, tmp_var);
      cmp175463_322 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_350_inst
    process(tmp495_345) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp495_345, type_cast_349_wire_constant, tmp_var);
      tmp496_351 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_567_inst
    process(tmp482_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp482_562, type_cast_566_wire_constant, tmp_var);
      tmp483_568 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1045_inst
    process(conv266_1037, conv268_781) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv266_1037, conv268_781, tmp_var);
      cmp269_1046 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_852_inst
    process(conv241_848, conv243_775) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv241_848, conv243_775, tmp_var);
      cmp244_853 <= tmp_var; --
    end process;
    -- shared split operator group (122) : array_obj_ref_1079_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom273_1078_scaled;
      array_obj_ref_1079_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1079_index_offset_req_0;
      array_obj_ref_1079_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1079_index_offset_req_1;
      array_obj_ref_1079_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_1102_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom277_1101_scaled;
      array_obj_ref_1102_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1102_index_offset_req_0;
      array_obj_ref_1102_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1102_index_offset_req_1;
      array_obj_ref_1102_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_1538_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1537_scaled;
      array_obj_ref_1538_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1538_index_offset_req_0;
      array_obj_ref_1538_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1538_index_offset_req_1;
      array_obj_ref_1538_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_389_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar489_388_scaled;
      array_obj_ref_389_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_389_index_offset_req_0;
      array_obj_ref_389_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_389_index_offset_req_1;
      array_obj_ref_389_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- shared split operator group (126) : array_obj_ref_606_index_offset 
    ApIntAdd_group_126: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_605_scaled;
      array_obj_ref_606_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_606_index_offset_req_0;
      array_obj_ref_606_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_606_index_offset_req_1;
      array_obj_ref_606_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_126_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_126_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_126",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 126
    -- shared split operator group (127) : array_obj_ref_876_index_offset 
    ApIntAdd_group_127: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom247_875_scaled;
      array_obj_ref_876_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_876_index_offset_req_0;
      array_obj_ref_876_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_876_index_offset_req_1;
      array_obj_ref_876_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_127_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_127_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_127",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 127
    -- shared split operator group (128) : array_obj_ref_899_index_offset 
    ApIntAdd_group_128: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom251_898_scaled;
      array_obj_ref_899_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_899_index_offset_req_0;
      array_obj_ref_899_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_899_index_offset_req_1;
      array_obj_ref_899_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_128_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_128_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_128",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 128
    -- unary operator type_cast_1367_inst
    process(call233_768) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call233_768, tmp_var);
      type_cast_1367_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1375_inst
    process(call310_1372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call310_1372, tmp_var);
      type_cast_1375_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1088_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1088_load_0_req_0;
      ptr_deref_1088_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1088_load_0_req_1;
      ptr_deref_1088_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen271_exec_guard_1025_delayed_7_0_1084(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1088_word_address_0;
      ptr_deref_1088_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1543_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1543_load_0_req_0;
      ptr_deref_1543_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1543_load_0_req_1;
      ptr_deref_1543_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1543_word_address_0;
      ptr_deref_1543_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_885_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_885_load_0_req_0;
      ptr_deref_885_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_885_load_0_req_1;
      ptr_deref_885_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen_exec_guard_876_delayed_7_0_881(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_885_word_address_0;
      ptr_deref_885_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : ptr_deref_1113_store_0 ptr_deref_910_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1113_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_910_store_0_req_0;
      ptr_deref_1113_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_910_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1113_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_910_store_0_req_1;
      ptr_deref_1113_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_910_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xthen_exec_guard_893_delayed_13_0_904(0);
      guard_vector(1)  <= ifx_xthen271_exec_guard_1042_delayed_13_0_1107(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1113_word_address_0 & ptr_deref_910_word_address_0;
      data_in <= ptr_deref_1113_data_0 & ptr_deref_910_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_526_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_526_store_0_req_0;
      ptr_deref_526_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_526_store_0_req_1;
      ptr_deref_526_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_526_word_address_0;
      data_in <= ptr_deref_526_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_743_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_743_store_0_req_0;
      ptr_deref_743_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_743_store_0_req_1;
      ptr_deref_743_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_743_word_address_0;
      data_in <= ptr_deref_743_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Concat_input_pipe_189_inst RPIPE_Concat_input_pipe_114_inst RPIPE_Concat_input_pipe_64_inst RPIPE_Concat_input_pipe_214_inst RPIPE_Concat_input_pipe_226_inst RPIPE_Concat_input_pipe_51_inst RPIPE_Concat_input_pipe_139_inst RPIPE_Concat_input_pipe_201_inst RPIPE_Concat_input_pipe_101_inst RPIPE_Concat_input_pipe_176_inst RPIPE_Concat_input_pipe_126_inst RPIPE_Concat_input_pipe_164_inst RPIPE_Concat_input_pipe_89_inst RPIPE_Concat_input_pipe_151_inst RPIPE_Concat_input_pipe_39_inst RPIPE_Concat_input_pipe_25_inst RPIPE_Concat_input_pipe_76_inst RPIPE_Concat_input_pipe_239_inst RPIPE_Concat_input_pipe_393_inst RPIPE_Concat_input_pipe_406_inst RPIPE_Concat_input_pipe_424_inst RPIPE_Concat_input_pipe_442_inst RPIPE_Concat_input_pipe_460_inst RPIPE_Concat_input_pipe_478_inst RPIPE_Concat_input_pipe_496_inst RPIPE_Concat_input_pipe_514_inst RPIPE_Concat_input_pipe_610_inst RPIPE_Concat_input_pipe_623_inst RPIPE_Concat_input_pipe_641_inst RPIPE_Concat_input_pipe_659_inst RPIPE_Concat_input_pipe_677_inst RPIPE_Concat_input_pipe_695_inst RPIPE_Concat_input_pipe_713_inst RPIPE_Concat_input_pipe_731_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_Concat_input_pipe_189_inst_req_0;
      reqL_unguarded(32) <= RPIPE_Concat_input_pipe_114_inst_req_0;
      reqL_unguarded(31) <= RPIPE_Concat_input_pipe_64_inst_req_0;
      reqL_unguarded(30) <= RPIPE_Concat_input_pipe_214_inst_req_0;
      reqL_unguarded(29) <= RPIPE_Concat_input_pipe_226_inst_req_0;
      reqL_unguarded(28) <= RPIPE_Concat_input_pipe_51_inst_req_0;
      reqL_unguarded(27) <= RPIPE_Concat_input_pipe_139_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Concat_input_pipe_201_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Concat_input_pipe_101_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Concat_input_pipe_176_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Concat_input_pipe_126_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Concat_input_pipe_164_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Concat_input_pipe_89_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Concat_input_pipe_151_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Concat_input_pipe_39_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Concat_input_pipe_25_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Concat_input_pipe_76_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Concat_input_pipe_239_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Concat_input_pipe_393_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Concat_input_pipe_406_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Concat_input_pipe_424_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Concat_input_pipe_442_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Concat_input_pipe_460_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Concat_input_pipe_478_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Concat_input_pipe_496_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Concat_input_pipe_514_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Concat_input_pipe_610_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Concat_input_pipe_623_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Concat_input_pipe_641_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Concat_input_pipe_659_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Concat_input_pipe_677_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Concat_input_pipe_695_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Concat_input_pipe_713_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Concat_input_pipe_731_inst_req_0;
      RPIPE_Concat_input_pipe_189_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_Concat_input_pipe_114_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_Concat_input_pipe_64_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_Concat_input_pipe_214_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_Concat_input_pipe_226_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_Concat_input_pipe_51_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_Concat_input_pipe_139_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Concat_input_pipe_201_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Concat_input_pipe_101_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Concat_input_pipe_176_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Concat_input_pipe_126_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Concat_input_pipe_164_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Concat_input_pipe_89_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Concat_input_pipe_151_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Concat_input_pipe_39_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Concat_input_pipe_25_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Concat_input_pipe_76_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Concat_input_pipe_239_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Concat_input_pipe_393_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Concat_input_pipe_406_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Concat_input_pipe_424_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Concat_input_pipe_442_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Concat_input_pipe_460_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Concat_input_pipe_478_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Concat_input_pipe_496_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Concat_input_pipe_514_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Concat_input_pipe_610_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Concat_input_pipe_623_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Concat_input_pipe_641_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Concat_input_pipe_659_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Concat_input_pipe_677_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Concat_input_pipe_695_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Concat_input_pipe_713_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Concat_input_pipe_731_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_Concat_input_pipe_189_inst_req_1;
      reqR_unguarded(32) <= RPIPE_Concat_input_pipe_114_inst_req_1;
      reqR_unguarded(31) <= RPIPE_Concat_input_pipe_64_inst_req_1;
      reqR_unguarded(30) <= RPIPE_Concat_input_pipe_214_inst_req_1;
      reqR_unguarded(29) <= RPIPE_Concat_input_pipe_226_inst_req_1;
      reqR_unguarded(28) <= RPIPE_Concat_input_pipe_51_inst_req_1;
      reqR_unguarded(27) <= RPIPE_Concat_input_pipe_139_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Concat_input_pipe_201_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Concat_input_pipe_101_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Concat_input_pipe_176_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Concat_input_pipe_126_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Concat_input_pipe_164_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Concat_input_pipe_89_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Concat_input_pipe_151_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Concat_input_pipe_39_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Concat_input_pipe_25_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Concat_input_pipe_76_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Concat_input_pipe_239_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Concat_input_pipe_393_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Concat_input_pipe_406_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Concat_input_pipe_424_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Concat_input_pipe_442_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Concat_input_pipe_460_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Concat_input_pipe_478_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Concat_input_pipe_496_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Concat_input_pipe_514_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Concat_input_pipe_610_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Concat_input_pipe_623_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Concat_input_pipe_641_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Concat_input_pipe_659_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Concat_input_pipe_677_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Concat_input_pipe_695_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Concat_input_pipe_713_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Concat_input_pipe_731_inst_req_1;
      RPIPE_Concat_input_pipe_189_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_Concat_input_pipe_114_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_Concat_input_pipe_64_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_Concat_input_pipe_214_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_Concat_input_pipe_226_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_Concat_input_pipe_51_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_Concat_input_pipe_139_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Concat_input_pipe_201_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Concat_input_pipe_101_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Concat_input_pipe_176_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Concat_input_pipe_126_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Concat_input_pipe_164_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Concat_input_pipe_89_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Concat_input_pipe_151_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Concat_input_pipe_39_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Concat_input_pipe_25_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Concat_input_pipe_76_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Concat_input_pipe_239_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Concat_input_pipe_393_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Concat_input_pipe_406_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Concat_input_pipe_424_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Concat_input_pipe_442_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Concat_input_pipe_460_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Concat_input_pipe_478_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Concat_input_pipe_496_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Concat_input_pipe_514_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Concat_input_pipe_610_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Concat_input_pipe_623_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Concat_input_pipe_641_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Concat_input_pipe_659_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Concat_input_pipe_677_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Concat_input_pipe_695_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Concat_input_pipe_713_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Concat_input_pipe_731_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call55_190 <= data_out(271 downto 264);
      call28_115 <= data_out(263 downto 256);
      call10_65 <= data_out(255 downto 248);
      call64_215 <= data_out(247 downto 240);
      call68_227 <= data_out(239 downto 232);
      call5_52 <= data_out(231 downto 224);
      call37_140 <= data_out(223 downto 216);
      call59_202 <= data_out(215 downto 208);
      call23_102 <= data_out(207 downto 200);
      call50_177 <= data_out(199 downto 192);
      call32_127 <= data_out(191 downto 184);
      call46_165 <= data_out(183 downto 176);
      call19_90 <= data_out(175 downto 168);
      call41_152 <= data_out(167 downto 160);
      call2_40 <= data_out(159 downto 152);
      call_26 <= data_out(151 downto 144);
      call14_77 <= data_out(143 downto 136);
      call73_240 <= data_out(135 downto 128);
      call124_394 <= data_out(127 downto 120);
      call128_407 <= data_out(119 downto 112);
      call134_425 <= data_out(111 downto 104);
      call140_443 <= data_out(103 downto 96);
      call146_461 <= data_out(95 downto 88);
      call152_479 <= data_out(87 downto 80);
      call158_497 <= data_out(79 downto 72);
      call164_515 <= data_out(71 downto 64);
      call180_611 <= data_out(63 downto 56);
      call184_624 <= data_out(55 downto 48);
      call190_642 <= data_out(47 downto 40);
      call196_660 <= data_out(39 downto 32);
      call202_678 <= data_out(31 downto 24);
      call208_696 <= data_out(23 downto 16);
      call214_714 <= data_out(15 downto 8);
      call220_732 <= data_out(7 downto 0);
      Concat_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Concat_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Concat_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Concat_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Concat_input_pipe_pipe_read_req(0),
          oack => Concat_input_pipe_pipe_read_ack(0),
          odata => Concat_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Concat_output_pipe_1457_inst WPIPE_Concat_output_pipe_1460_inst WPIPE_Concat_output_pipe_1463_inst WPIPE_Concat_output_pipe_1466_inst WPIPE_Concat_output_pipe_1469_inst WPIPE_Concat_output_pipe_1472_inst WPIPE_Concat_output_pipe_1475_inst WPIPE_Concat_output_pipe_1478_inst WPIPE_Concat_output_pipe_1619_inst WPIPE_Concat_output_pipe_1622_inst WPIPE_Concat_output_pipe_1625_inst WPIPE_Concat_output_pipe_1628_inst WPIPE_Concat_output_pipe_1631_inst WPIPE_Concat_output_pipe_1634_inst WPIPE_Concat_output_pipe_1637_inst WPIPE_Concat_output_pipe_1640_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Concat_output_pipe_1457_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Concat_output_pipe_1460_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Concat_output_pipe_1463_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Concat_output_pipe_1466_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Concat_output_pipe_1469_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Concat_output_pipe_1472_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Concat_output_pipe_1475_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Concat_output_pipe_1478_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Concat_output_pipe_1619_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Concat_output_pipe_1622_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Concat_output_pipe_1625_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Concat_output_pipe_1628_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Concat_output_pipe_1631_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Concat_output_pipe_1634_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Concat_output_pipe_1637_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Concat_output_pipe_1640_inst_req_0;
      WPIPE_Concat_output_pipe_1457_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1460_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1463_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1466_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1469_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1472_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1475_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1478_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1619_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1622_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1625_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1628_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1631_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1634_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1637_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1640_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Concat_output_pipe_1457_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Concat_output_pipe_1460_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Concat_output_pipe_1463_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Concat_output_pipe_1466_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Concat_output_pipe_1469_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Concat_output_pipe_1472_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Concat_output_pipe_1475_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Concat_output_pipe_1478_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Concat_output_pipe_1619_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Concat_output_pipe_1622_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Concat_output_pipe_1625_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Concat_output_pipe_1628_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Concat_output_pipe_1631_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Concat_output_pipe_1634_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Concat_output_pipe_1637_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Concat_output_pipe_1640_inst_req_1;
      WPIPE_Concat_output_pipe_1457_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1460_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1463_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1466_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1469_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1472_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1475_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1478_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1619_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1622_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1625_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1628_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1631_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1634_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1637_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1640_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv359_1456 & conv353_1446 & conv347_1436 & conv341_1426 & conv335_1416 & conv329_1406 & conv323_1396 & conv317_1386 & conv435_1618 & conv429_1608 & conv423_1598 & conv417_1588 & conv411_1578 & conv405_1568 & conv399_1558 & conv393_1548;
      Concat_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Concat_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Concat_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Concat_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Concat_output_pipe_pipe_write_req(0),
          oack => Concat_output_pipe_pipe_write_ack(0),
          odata => Concat_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_768_call call_stmt_1372_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_768_call_req_0;
      reqL_unguarded(0) <= call_stmt_1372_call_req_0;
      call_stmt_768_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1372_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_768_call_req_1;
      reqR_unguarded(0) <= call_stmt_1372_call_req_1;
      call_stmt_768_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1372_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call233_768 <= data_out(127 downto 64);
      call310_1372 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end concat_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_14_inst_req_0 : boolean;
  signal WPIPE_timer_req_14_inst_ack_0 : boolean;
  signal WPIPE_timer_req_14_inst_req_1 : boolean;
  signal WPIPE_timer_req_14_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_19_inst_req_0 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_19_inst_req_1 : boolean;
  signal RPIPE_timer_resp_19_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/req
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_start_
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_19_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_14_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_sample_completed_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_start_
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Sample/ack
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$entry
      -- CP-element group 1: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_14_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_update_completed_
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/$exit
      -- CP-element group 2: 	 assign_stmt_17_to_assign_stmt_20/WPIPE_timer_req_14_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_14_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_start_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_sample_completed_
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Sample/ra
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$entry
      -- CP-element group 3: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_19_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_update_completed_
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/$exit
      -- CP-element group 4: 	 assign_stmt_17_to_assign_stmt_20/RPIPE_timer_resp_19_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_19_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_17_to_assign_stmt_20/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_16_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_16_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_19_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_19_inst_req_0;
      RPIPE_timer_resp_19_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_19_inst_req_1;
      RPIPE_timer_resp_19_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_14_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_0;
      WPIPE_timer_req_14_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_14_inst_req_1;
      WPIPE_timer_req_14_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_16_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3761_start: Boolean;
  signal timerDaemon_CP_3761_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1677_branch_req_0 : boolean;
  signal RPIPE_timer_req_1686_inst_ack_1 : boolean;
  signal phi_stmt_1679_ack_0 : boolean;
  signal phi_stmt_1679_req_1 : boolean;
  signal nCOUNTER_1692_1683_buf_req_0 : boolean;
  signal nCOUNTER_1692_1683_buf_ack_0 : boolean;
  signal phi_stmt_1679_req_0 : boolean;
  signal RPIPE_timer_req_1686_inst_ack_0 : boolean;
  signal RPIPE_timer_req_1686_inst_req_0 : boolean;
  signal RPIPE_timer_req_1686_inst_req_1 : boolean;
  signal nCOUNTER_1692_1683_buf_req_1 : boolean;
  signal nCOUNTER_1692_1683_buf_ack_1 : boolean;
  signal WPIPE_timer_resp_1694_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1694_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_1694_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1694_inst_ack_1 : boolean;
  signal do_while_stmt_1677_branch_ack_0 : boolean;
  signal do_while_stmt_1677_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3761_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3761_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3761_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3761_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3761: Block -- control-path 
    signal timerDaemon_CP_3761_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3761_elements(0) <= timerDaemon_CP_3761_start;
    timerDaemon_CP_3761_symbol <= timerDaemon_CP_3761_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1676/branch_block_stmt_1676__entry__
      -- CP-element group 0: 	 branch_block_stmt_1676/do_while_stmt_1677__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1676/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1676/branch_block_stmt_1676__exit__
      -- CP-element group 1: 	 branch_block_stmt_1676/do_while_stmt_1677__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1676/$exit
      -- 
    timerDaemon_CP_3761_elements(1) <= timerDaemon_CP_3761_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677__entry__
      -- CP-element group 2: 	 branch_block_stmt_1676/do_while_stmt_1677/$entry
      -- 
    timerDaemon_CP_3761_elements(2) <= timerDaemon_CP_3761_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677__exit__
      -- 
    -- Element group timerDaemon_CP_3761_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_back
      -- 
    -- Element group timerDaemon_CP_3761_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/$entry
      -- 
    timerDaemon_CP_3761_elements(5) <= timerDaemon_CP_3761_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_body_done
      -- 
    timerDaemon_CP_3761_elements(6) <= timerDaemon_CP_3761_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3761_elements(7) <= timerDaemon_CP_3761_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3761_elements(8) <= timerDaemon_CP_3761_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_sample_start_
      -- 
    -- Element group timerDaemon_CP_3761_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/condition_evaluated
      -- 
    condition_evaluated_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(10), ack => do_while_stmt_1677_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(14) & timerDaemon_CP_3761_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(9) & timerDaemon_CP_3761_elements(15) & timerDaemon_CP_3761_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(17) & timerDaemon_CP_3761_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(16) & timerDaemon_CP_3761_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(18) & timerDaemon_CP_3761_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(9) & timerDaemon_CP_3761_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(9) & timerDaemon_CP_3761_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_3761_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_3761_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_trigger
      -- 
    timerDaemon_CP_3761_elements(19) <= timerDaemon_CP_3761_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_loopback_sample_req_ps
      -- 
    phi_stmt_1679_loopback_sample_req_3800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1679_loopback_sample_req_3800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(20), ack => phi_stmt_1679_req_1); -- 
    -- Element group timerDaemon_CP_3761_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_trigger
      -- 
    timerDaemon_CP_3761_elements(21) <= timerDaemon_CP_3761_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_entry_sample_req_ps
      -- 
    phi_stmt_1679_entry_sample_req_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1679_entry_sample_req_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(22), ack => phi_stmt_1679_req_0); -- 
    -- Element group timerDaemon_CP_3761_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1679_phi_mux_ack_ps
      -- 
    phi_stmt_1679_phi_mux_ack_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1679_ack_0, ack => timerDaemon_CP_3761_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_3761_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_start__ps
      -- 
    -- Element group timerDaemon_CP_3761_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_completed__ps
      -- 
    timerDaemon_CP_3761_elements(26) <= timerDaemon_CP_3761_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/type_cast_1682_update_completed_
      -- 
    -- Element group timerDaemon_CP_3761_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_3761_elements(25), ack => timerDaemon_CP_3761_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/req
      -- 
    req_3827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(28), ack => nCOUNTER_1692_1683_buf_req_0); -- 
    -- Element group timerDaemon_CP_3761_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/$entry
      -- 
    req_3832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(29), ack => nCOUNTER_1692_1683_buf_req_1); -- 
    -- Element group timerDaemon_CP_3761_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_sample_completed__ps
      -- 
    ack_3828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1692_1683_buf_ack_0, ack => timerDaemon_CP_3761_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/R_nCOUNTER_1683_update_completed__ps
      -- 
    ack_3833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1692_1683_buf_ack_1, ack => timerDaemon_CP_3761_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(9) & timerDaemon_CP_3761_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/rr
      -- 
    rr_3846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(33), ack => RPIPE_timer_req_1686_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(11) & timerDaemon_CP_3761_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/$entry
      -- 
    cr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(34), ack => RPIPE_timer_req_1686_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(13) & timerDaemon_CP_3761_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Sample/$exit
      -- 
    ra_3847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1686_inst_ack_0, ack => timerDaemon_CP_3761_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/phi_stmt_1684_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/RPIPE_timer_req_1686_Update/$exit
      -- 
    ca_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1686_inst_ack_1, ack => timerDaemon_CP_3761_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/req
      -- 
    req_3860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(37), ack => WPIPE_timer_resp_1694_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(18) & timerDaemon_CP_3761_elements(36) & timerDaemon_CP_3761_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/req
      -- 
    ack_3861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1694_inst_ack_0, ack => timerDaemon_CP_3761_elements(38)); -- 
    req_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3761_elements(38), ack => WPIPE_timer_resp_1694_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/WPIPE_timer_resp_1694_Update/ack
      -- 
    ack_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1694_inst_ack_1, ack => timerDaemon_CP_3761_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3761_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_3761_elements(9), ack => timerDaemon_CP_3761_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1676/do_while_stmt_1677/do_while_stmt_1677_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3761_elements(12) & timerDaemon_CP_3761_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3761_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_exit/ack
      -- 
    ack_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1677_branch_ack_0, ack => timerDaemon_CP_3761_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1676/do_while_stmt_1677/loop_taken/ack
      -- 
    ack_3875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1677_branch_ack_1, ack => timerDaemon_CP_3761_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1676/do_while_stmt_1677/$exit
      -- 
    timerDaemon_CP_3761_elements(44) <= timerDaemon_CP_3761_elements(3);
    timerDaemon_do_while_stmt_1677_terminator_3876: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1677_terminator_3876", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_3761_elements(6),loop_continue => timerDaemon_CP_3761_elements(43),loop_terminate => timerDaemon_CP_3761_elements(42),loop_back => timerDaemon_CP_3761_elements(4),loop_exit => timerDaemon_CP_3761_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1679_phi_seq_3834_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3761_elements(21);
      timerDaemon_CP_3761_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3761_elements(24);
      timerDaemon_CP_3761_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3761_elements(26);
      timerDaemon_CP_3761_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3761_elements(19);
      timerDaemon_CP_3761_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3761_elements(30);
      timerDaemon_CP_3761_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3761_elements(31);
      timerDaemon_CP_3761_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1679_phi_seq_3834 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1679_phi_seq_3834") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3761_elements(11), 
          phi_sample_ack => timerDaemon_CP_3761_elements(17), 
          phi_update_req => timerDaemon_CP_3761_elements(13), 
          phi_update_ack => timerDaemon_CP_3761_elements(18), 
          phi_mux_ack => timerDaemon_CP_3761_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3786_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3761_elements(7);
        preds(1)  <= timerDaemon_CP_3761_elements(8);
        entry_tmerge_3786 : transition_merge -- 
          generic map(name => " entry_tmerge_3786")
          port map (preds => preds, symbol_out => timerDaemon_CP_3761_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1679 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1686_wire : std_logic_vector(0 downto 0);
    signal konst_1690_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1698_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1692 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1692_1683_buffered : std_logic_vector(63 downto 0);
    signal req_1684 : std_logic_vector(0 downto 0);
    signal type_cast_1682_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1690_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1698_wire_constant <= "1";
    type_cast_1682_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1679: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1682_wire_constant & nCOUNTER_1692_1683_buffered;
      req <= phi_stmt_1679_req_0 & phi_stmt_1679_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1679",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1679_ack_0,
          idata => idata,
          odata => COUNTER_1679,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1679
    nCOUNTER_1692_1683_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1692_1683_buf_req_0;
      nCOUNTER_1692_1683_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1692_1683_buf_req_1;
      nCOUNTER_1692_1683_buf_ack_1<= rack(0);
      nCOUNTER_1692_1683_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1692_1683_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1692_1683_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1684
    process(RPIPE_timer_req_1686_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1686_wire(0 downto 0);
      req_1684 <= tmp_var; -- 
    end process;
    do_while_stmt_1677_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1698_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1677_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1677_branch_req_0,
          ack0 => do_while_stmt_1677_branch_ack_0,
          ack1 => do_while_stmt_1677_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1691_inst
    process(COUNTER_1679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1679, konst_1690_wire_constant, tmp_var);
      nCOUNTER_1692 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1686_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1686_inst_req_0;
      RPIPE_timer_req_1686_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1686_inst_req_1;
      RPIPE_timer_req_1686_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1686_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1694_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1694_inst_req_0;
      WPIPE_timer_resp_1694_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1694_inst_req_1;
      WPIPE_timer_resp_1694_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1684(0);
      data_in <= COUNTER_1679;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Concat_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Concat_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module concat
  component concat is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module concat
  signal concat_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal concat_tag_out   : std_logic_vector(1 downto 0);
  signal concat_start_req : std_logic;
  signal concat_start_ack : std_logic;
  signal concat_fin_req   : std_logic;
  signal concat_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe Concat_input_pipe
  signal Concat_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal Concat_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal Concat_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Concat_output_pipe
  signal Concat_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Concat_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Concat_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module concat
  concat_instance:concat-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => concat_start_req,
      start_ack => concat_start_ack,
      fin_req => concat_fin_req,
      fin_ack => concat_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      Concat_input_pipe_pipe_read_req => Concat_input_pipe_pipe_read_req(0 downto 0),
      Concat_input_pipe_pipe_read_ack => Concat_input_pipe_pipe_read_ack(0 downto 0),
      Concat_input_pipe_pipe_read_data => Concat_input_pipe_pipe_read_data(7 downto 0),
      Concat_output_pipe_pipe_write_req => Concat_output_pipe_pipe_write_req(0 downto 0),
      Concat_output_pipe_pipe_write_ack => Concat_output_pipe_pipe_write_ack(0 downto 0),
      Concat_output_pipe_pipe_write_data => Concat_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => concat_tag_in,
      tag_out => concat_tag_out-- 
    ); -- 
  -- module will be run forever 
  concat_tag_in <= (others => '0');
  concat_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => concat_start_req, start_ack => concat_start_ack,  fin_req => concat_fin_req,  fin_ack => concat_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  Concat_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_input_pipe_pipe_read_req,
      read_ack => Concat_input_pipe_pipe_read_ack,
      read_data => Concat_input_pipe_pipe_read_data,
      write_req => Concat_input_pipe_pipe_write_req,
      write_ack => Concat_input_pipe_pipe_write_ack,
      write_data => Concat_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Concat_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_output_pipe_pipe_read_req,
      read_ack => Concat_output_pipe_pipe_read_ack,
      read_data => Concat_output_pipe_pipe_read_data,
      write_req => Concat_output_pipe_pipe_write_req,
      write_ack => Concat_output_pipe_pipe_write_ack,
      write_data => Concat_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
