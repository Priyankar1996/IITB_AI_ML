-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_727_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_1 : boolean;
  signal if_stmt_632_branch_ack_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal addr_of_689_final_reg_ack_1 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_1332_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal type_cast_1048_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_1 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal if_stmt_632_branch_req_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_req_1 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_1 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_1 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_req_1 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_ack_0 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_0 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_0 : boolean;
  signal type_cast_339_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_1 : boolean;
  signal type_cast_339_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_1 : boolean;
  signal type_cast_696_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_0 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal array_obj_ref_688_index_offset_req_0 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_1048_inst_ack_0 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_0 : boolean;
  signal type_cast_696_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_req_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_1 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_1 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal type_cast_556_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_1 : boolean;
  signal type_cast_1048_inst_req_1 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal type_cast_556_inst_req_1 : boolean;
  signal type_cast_259_inst_req_0 : boolean;
  signal type_cast_259_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_0 : boolean;
  signal type_cast_259_inst_req_1 : boolean;
  signal type_cast_259_inst_ack_1 : boolean;
  signal type_cast_556_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_0 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal type_cast_556_inst_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_1048_inst_ack_1 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 : boolean;
  signal type_cast_289_inst_req_0 : boolean;
  signal type_cast_289_inst_ack_0 : boolean;
  signal type_cast_289_inst_req_1 : boolean;
  signal type_cast_289_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_314_inst_req_0 : boolean;
  signal type_cast_314_inst_ack_0 : boolean;
  signal type_cast_314_inst_req_1 : boolean;
  signal type_cast_314_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_0 : boolean;
  signal if_stmt_632_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 : boolean;
  signal type_cast_327_inst_req_0 : boolean;
  signal type_cast_327_inst_ack_0 : boolean;
  signal type_cast_327_inst_req_1 : boolean;
  signal type_cast_327_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 : boolean;
  signal type_cast_352_inst_req_0 : boolean;
  signal type_cast_352_inst_ack_0 : boolean;
  signal type_cast_352_inst_req_1 : boolean;
  signal type_cast_352_inst_ack_1 : boolean;
  signal type_cast_1400_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal type_cast_364_inst_req_0 : boolean;
  signal type_cast_364_inst_ack_0 : boolean;
  signal type_cast_364_inst_req_1 : boolean;
  signal type_cast_364_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal type_cast_377_inst_req_0 : boolean;
  signal type_cast_377_inst_ack_0 : boolean;
  signal type_cast_377_inst_req_1 : boolean;
  signal type_cast_377_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_1 : boolean;
  signal type_cast_389_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_0 : boolean;
  signal type_cast_389_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal type_cast_402_inst_req_0 : boolean;
  signal type_cast_402_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 : boolean;
  signal type_cast_402_inst_req_1 : boolean;
  signal type_cast_402_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_0 : boolean;
  signal type_cast_1332_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal if_stmt_416_branch_req_0 : boolean;
  signal if_stmt_416_branch_ack_1 : boolean;
  signal if_stmt_416_branch_ack_0 : boolean;
  signal if_stmt_431_branch_req_0 : boolean;
  signal if_stmt_431_branch_ack_1 : boolean;
  signal if_stmt_431_branch_ack_0 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal array_obj_ref_481_index_offset_req_0 : boolean;
  signal array_obj_ref_481_index_offset_ack_0 : boolean;
  signal array_obj_ref_481_index_offset_req_1 : boolean;
  signal array_obj_ref_481_index_offset_ack_1 : boolean;
  signal addr_of_482_final_reg_req_0 : boolean;
  signal addr_of_482_final_reg_ack_0 : boolean;
  signal addr_of_482_final_reg_req_1 : boolean;
  signal addr_of_482_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 : boolean;
  signal type_cast_489_inst_req_0 : boolean;
  signal type_cast_489_inst_ack_0 : boolean;
  signal type_cast_489_inst_req_1 : boolean;
  signal type_cast_489_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 : boolean;
  signal type_cast_502_inst_req_0 : boolean;
  signal type_cast_502_inst_ack_0 : boolean;
  signal type_cast_502_inst_req_1 : boolean;
  signal type_cast_502_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_1 : boolean;
  signal type_cast_745_inst_req_0 : boolean;
  signal type_cast_745_inst_ack_0 : boolean;
  signal type_cast_745_inst_req_1 : boolean;
  signal type_cast_745_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal type_cast_1400_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_0 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_1 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 : boolean;
  signal type_cast_1370_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_0 : boolean;
  signal type_cast_1400_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 : boolean;
  signal type_cast_1370_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_0 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_0 : boolean;
  signal ptr_deref_825_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_0 : boolean;
  signal ptr_deref_825_store_0_ack_0 : boolean;
  signal ptr_deref_825_store_0_req_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_0 : boolean;
  signal ptr_deref_825_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_1 : boolean;
  signal type_cast_1400_inst_req_0 : boolean;
  signal if_stmt_839_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal if_stmt_839_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal if_stmt_839_branch_ack_0 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal type_cast_850_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal type_cast_850_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_1 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_858_inst_req_0 : boolean;
  signal type_cast_858_inst_ack_0 : boolean;
  signal type_cast_858_inst_req_1 : boolean;
  signal type_cast_858_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 : boolean;
  signal if_stmt_876_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal if_stmt_876_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal if_stmt_876_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_0 : boolean;
  signal array_obj_ref_932_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal array_obj_ref_932_index_offset_ack_0 : boolean;
  signal array_obj_ref_932_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal array_obj_ref_932_index_offset_ack_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_0 : boolean;
  signal addr_of_933_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal addr_of_933_final_reg_ack_0 : boolean;
  signal ptr_deref_1366_load_0_req_0 : boolean;
  signal addr_of_933_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal addr_of_933_final_reg_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal ptr_deref_936_store_0_req_0 : boolean;
  signal ptr_deref_936_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal ptr_deref_936_store_0_req_1 : boolean;
  signal ptr_deref_936_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_1 : boolean;
  signal type_cast_1420_inst_req_0 : boolean;
  signal if_stmt_951_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_0 : boolean;
  signal if_stmt_951_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal if_stmt_951_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_1 : boolean;
  signal call_stmt_962_call_req_0 : boolean;
  signal call_stmt_962_call_ack_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_1 : boolean;
  signal call_stmt_962_call_req_1 : boolean;
  signal call_stmt_962_call_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_972_inst_req_0 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_969_inst_req_0 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_969_inst_req_1 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_1 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal type_cast_1370_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_1 : boolean;
  signal type_cast_1370_inst_req_0 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1410_inst_ack_1 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1106_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1106_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1106_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1106_inst_ack_1 : boolean;
  signal type_cast_1410_inst_req_1 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 : boolean;
  signal type_cast_1390_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_0 : boolean;
  signal type_cast_1390_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_1 : boolean;
  signal if_stmt_1305_branch_ack_0 : boolean;
  signal ptr_deref_1366_load_0_ack_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_1 : boolean;
  signal ptr_deref_1366_load_0_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_0 : boolean;
  signal type_cast_1390_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal addr_of_1362_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal addr_of_1362_final_reg_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal if_stmt_1305_branch_ack_1 : boolean;
  signal type_cast_1390_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal addr_of_1362_final_reg_ack_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal addr_of_1362_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal type_cast_1440_inst_ack_1 : boolean;
  signal type_cast_1440_inst_req_1 : boolean;
  signal if_stmt_1305_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_0 : boolean;
  signal type_cast_1440_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_1 : boolean;
  signal type_cast_1440_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_1 : boolean;
  signal type_cast_1160_inst_req_0 : boolean;
  signal array_obj_ref_1361_index_offset_ack_1 : boolean;
  signal type_cast_1160_inst_ack_0 : boolean;
  signal type_cast_1410_inst_ack_0 : boolean;
  signal type_cast_1160_inst_req_1 : boolean;
  signal array_obj_ref_1361_index_offset_req_1 : boolean;
  signal type_cast_1160_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1162_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1162_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1162_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1162_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_1 : boolean;
  signal type_cast_1430_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 : boolean;
  signal type_cast_1430_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_0 : boolean;
  signal type_cast_1410_inst_req_0 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal array_obj_ref_1361_index_offset_ack_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal array_obj_ref_1361_index_offset_req_0 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal ptr_deref_1366_load_0_ack_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_0 : boolean;
  signal type_cast_1430_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_1 : boolean;
  signal type_cast_1430_inst_req_0 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal type_cast_1420_inst_ack_1 : boolean;
  signal type_cast_1420_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1182_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1182_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1182_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1182_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 : boolean;
  signal type_cast_1420_inst_ack_0 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1185_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1185_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1185_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1185_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1188_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1188_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1188_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1188_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1191_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1191_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1191_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1191_inst_ack_1 : boolean;
  signal call_stmt_1195_call_req_0 : boolean;
  signal call_stmt_1195_call_ack_0 : boolean;
  signal call_stmt_1195_call_req_1 : boolean;
  signal call_stmt_1195_call_ack_1 : boolean;
  signal type_cast_1199_inst_req_0 : boolean;
  signal type_cast_1199_inst_ack_0 : boolean;
  signal type_cast_1199_inst_req_1 : boolean;
  signal type_cast_1199_inst_ack_1 : boolean;
  signal type_cast_1208_inst_req_0 : boolean;
  signal type_cast_1208_inst_ack_0 : boolean;
  signal type_cast_1208_inst_req_1 : boolean;
  signal type_cast_1208_inst_ack_1 : boolean;
  signal type_cast_1218_inst_req_0 : boolean;
  signal type_cast_1218_inst_ack_0 : boolean;
  signal type_cast_1218_inst_req_1 : boolean;
  signal type_cast_1218_inst_ack_1 : boolean;
  signal type_cast_1228_inst_req_0 : boolean;
  signal type_cast_1228_inst_ack_0 : boolean;
  signal type_cast_1228_inst_req_1 : boolean;
  signal type_cast_1228_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_1248_inst_req_0 : boolean;
  signal type_cast_1248_inst_ack_0 : boolean;
  signal type_cast_1248_inst_req_1 : boolean;
  signal type_cast_1248_inst_ack_1 : boolean;
  signal type_cast_1258_inst_req_0 : boolean;
  signal type_cast_1258_inst_ack_0 : boolean;
  signal type_cast_1258_inst_req_1 : boolean;
  signal type_cast_1258_inst_ack_1 : boolean;
  signal type_cast_1268_inst_req_0 : boolean;
  signal type_cast_1268_inst_ack_0 : boolean;
  signal type_cast_1268_inst_req_1 : boolean;
  signal type_cast_1268_inst_ack_1 : boolean;
  signal type_cast_1278_inst_req_0 : boolean;
  signal type_cast_1278_inst_ack_0 : boolean;
  signal type_cast_1278_inst_req_1 : boolean;
  signal type_cast_1278_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1 : boolean;
  signal if_stmt_1477_branch_req_0 : boolean;
  signal if_stmt_1477_branch_ack_1 : boolean;
  signal if_stmt_1477_branch_ack_0 : boolean;
  signal phi_stmt_469_req_0 : boolean;
  signal type_cast_475_inst_req_0 : boolean;
  signal type_cast_475_inst_ack_0 : boolean;
  signal type_cast_475_inst_req_1 : boolean;
  signal type_cast_475_inst_ack_1 : boolean;
  signal phi_stmt_469_req_1 : boolean;
  signal phi_stmt_469_ack_0 : boolean;
  signal phi_stmt_676_req_1 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal phi_stmt_676_req_0 : boolean;
  signal phi_stmt_676_ack_0 : boolean;
  signal phi_stmt_920_req_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal phi_stmt_920_req_0 : boolean;
  signal phi_stmt_920_ack_0 : boolean;
  signal phi_stmt_1349_req_0 : boolean;
  signal type_cast_1355_inst_req_0 : boolean;
  signal type_cast_1355_inst_ack_0 : boolean;
  signal type_cast_1355_inst_req_1 : boolean;
  signal type_cast_1355_inst_ack_1 : boolean;
  signal phi_stmt_1349_req_1 : boolean;
  signal phi_stmt_1349_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(496 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(496);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_339_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_210_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_214_inst_req_1); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_255_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_259_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_263_inst_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_267_inst_req_1); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_289_inst_req_1); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_302_inst_req_1); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_314_inst_req_1); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_327_inst_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_352_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_364_inst_req_1); -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_377_inst_req_1); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_389_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_402_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_76_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_101_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_113_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_138_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_151_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_163_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_176_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_188_inst_req_0); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/rr
      -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_210_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/rr
      -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_214_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_218_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/rr
      -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_255_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/rr
      -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_259_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: 	44 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/rr
      -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_263_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(44);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/rr
      -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_267_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/ra
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/ca
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/cr
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/rr
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_289_inst_req_0); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/ra
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/ca
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/cr
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/rr
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_302_inst_req_0); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/ra
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_314_inst_req_0); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/ra
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/ca
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/cr
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/rr
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_327_inst_req_0); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/ra
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/ca
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/cr
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$entry
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_339_inst_req_0); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$exit
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_completed_
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/cr
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/rr
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_352_inst_req_0); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/cr
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/rr
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_364_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_377_inst_req_0); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/ra
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/cr
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/rr
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_389_inst_req_0); -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/ra
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/ca
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/cr
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/rr
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_402_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__exit__
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416__entry__
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_32/R_cmp513_417_place
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_else_link/$entry
      -- 
    branch_req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_416_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph515_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/dummy
      -- 
    if_choice_transition_908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_0); -- 
    cr_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	469 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	469 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/dummy
      -- 
    if_choice_transition_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_1); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	469 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	482 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/ra
      -- 
    ra_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	470 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__exit__
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- 
    ca_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	475 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/ack
      -- 
    ack_982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	475 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/req
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_482_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/ack
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	475 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/ack
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	475 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/cr
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/rr
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_489_inst_req_0); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/ra
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	475 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/cr
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/rr
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_502_inst_req_0); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/ra
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	475 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/ca
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_start_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_520_inst_req_0); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/ra
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	475 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/ca
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_start_
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_538_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_completed_
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	475 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$exit
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$exit
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$exit
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_556_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_completed_
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	475 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_completed_
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_completed_
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_completed_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_574_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_completed_
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	475 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_completed_
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_completed_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_start_
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_0); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_592_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_completed_
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	475 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/ca
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_completed_
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_completed_
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_610_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_completed_
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	475 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_completed_
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$entry
      -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_618_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$exit
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	475 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_completed_
      -- 
    ca_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__exit__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632__entry__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/R_exitcond3_633_place
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$exit
      -- 
    branch_req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_632_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	469 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	471 
    -- CP-element group 166: 	472 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_0); -- 
    cr_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_completed_
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	476 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__exit__
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	481 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_sample_complete
      -- 
    ack_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	481 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_ack
      -- 
    ack_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_689_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$exit
      -- 
    ack_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	481 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_ack
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	481 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_start_
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_696_inst_req_0); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	481 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_completed_
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_completed_
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_start_
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_709_inst_req_0); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$exit
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	481 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$exit
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_start_
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_start_
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_727_inst_req_0); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_completed_
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	481 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_completed_
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_start_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/ra
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/rr
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_745_inst_req_0); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/ra
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	481 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/ca
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_start_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/cr
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/rr
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_763_inst_req_0); -- 
    rr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/ra
      -- 
    ra_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	481 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/ca
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_start_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/cr
      -- 
    ra_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/rr
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_781_inst_req_0); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/ra
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	481 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/ca
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_start_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/cr
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/rr
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_799_inst_req_0); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/ra
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	481 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/ca
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_start_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/cr
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/rr
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_817_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/ra
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	481 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/ca
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/rr
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_825_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176) & convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	481 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/ca
      -- 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	169 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__exit__
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839__entry__
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_32/R_exitcond2_840_place
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_else_link/$entry
      -- 
    branch_req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_839_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(169) & convTranspose_CP_39_elements(207);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	482 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	477 
    -- CP-element group 210: 	478 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_0); -- 
    cr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	482 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	482 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/ca
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	482 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	482 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	482 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/ra
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	482 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__exit__
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876__entry__
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_32/R_cmp264505_877_place
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_else_link/$entry
      -- 
    branch_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_876_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__entry__
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph507_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/dummy
      -- 
    if_choice_transition_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_0); -- 
    cr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	489 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/ra
      -- 
    ra_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	483 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- 
    ca_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	488 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/ack
      -- 
    ack_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	488 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/req
      -- 
    ack_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_933_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	488 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/rr
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_936_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/ra
      -- 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	488 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__exit__
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951__entry__
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_32/R_exitcond_952_place
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_else_link/$entry
      -- 
    branch_req_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_951_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	489 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	484 
    -- CP-element group 230: 	485 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_0); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	489 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/cra
      -- 
    cra_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	489 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/rr
      -- 
    cca_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_967_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/ra
      -- 
    ra_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	489 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	373 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/ca
      -- 
    ca_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	489 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_969_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/$entry
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_972_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/req
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_update_start_
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_972_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_update_completed_
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/ack
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/req
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_sample_completed_
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_update_completed_
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/req
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_update_start_
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_sample_completed_
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/$entry
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/req
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_update_start_
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_update_completed_
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_update_start_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/req
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_996_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/req
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_sample_completed_
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_996_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_update_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_1000_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/ack
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_1000_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/$exit
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_1004_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/req
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_sample_completed_
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_1004_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_update_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_1007_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_sample_completed_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_1007_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_1010_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/req
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_1010_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	489 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/req
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_sample_completed_
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_1013_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/req
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_1016_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/req
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_update_start_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/$entry
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_1016_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_sample_start_
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/req
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_update_start_
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_update_completed_
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/req
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_update_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/req
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/$exit
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/req
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1034_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/req
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_update_start_
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_sample_completed_
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1034_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_update_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_sample_completed_
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_update_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	489 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/ra
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	489 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/ca
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/req
      -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1050_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/req
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_0, ack => convTranspose_CP_39_elements(284)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1050_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/ack
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_1, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	489 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_sample_completed_
      -- 
    ra_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	489 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_update_completed_
      -- 
    ca_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => convTranspose_CP_39_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_sample_start_
      -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1057_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(285) & convTranspose_CP_39_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1057_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_sample_start_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block1_start_1060_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/req
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_update_start_
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_sample_completed_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block1_start_1060_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/$entry
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block1_start_1063_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/req
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1063_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/$exit
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1066_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/req
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_sample_completed_
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block1_start_1066_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_update_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	489 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_update_start_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/req
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/$exit
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1069_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/$entry
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1072_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/req
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_update_start_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1072_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_update_completed_
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/$exit
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_sample_start_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_sample_completed_
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_update_completed_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_update_start_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/ack
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/$exit
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_update_start_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_sample_start_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/req
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/req
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block2_start_1090_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_update_start_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/req
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block2_start_1090_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/req
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block2_start_1093_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_update_start_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/req
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block2_start_1093_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/ack
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	489 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	489 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/req
      -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block2_start_1106_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_update_start_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1106_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block2_start_1106_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/ack
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1106_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	489 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	489 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/req
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1113_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_update_start_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1113_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1116_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_update_start_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1116_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	489 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_update_start_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block3_start_1125_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block3_start_1128_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_update_start_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block3_start_1128_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block3_start_1146_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_update_start_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block3_start_1146_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block3_start_1149_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_update_start_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block3_start_1149_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	489 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/ra
      -- 
    ra_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	489 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/ca
      -- 
    ca_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/req
      -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block3_start_1162_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(348) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_update_start_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1162_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block3_start_1162_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/ack
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1162_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	489 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/ra
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	489 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/ca
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/req
      -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block3_start_1169_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(353) & convTranspose_CP_39_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_update_start_
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block3_start_1169_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block3_start_1172_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_update_start_
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block3_start_1172_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_1, ack => convTranspose_CP_39_elements(360)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/ack
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	489 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_update_start_
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/cr
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1182_inst_ack_0, ack => convTranspose_CP_39_elements(365)); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => RPIPE_Block0_done_1182_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1182_inst_ack_1, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	489 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_update_start_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/cr
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1185_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => RPIPE_Block1_done_1185_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1185_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	489 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_update_start_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/cr
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1188_inst_ack_0, ack => convTranspose_CP_39_elements(369)); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => RPIPE_Block2_done_1188_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1188_inst_ack_1, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	489 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_update_start_
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/cr
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1191_inst_ack_0, ack => convTranspose_CP_39_elements(371)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => RPIPE_Block3_done_1191_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1191_inst_ack_1, ack => convTranspose_CP_39_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	234 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373: 	379 
    -- CP-element group 373: 	381 
    -- CP-element group 373: 	383 
    -- CP-element group 373: 	385 
    -- CP-element group 373: 	387 
    -- CP-element group 373: 	389 
    -- CP-element group 373: 	391 
    -- CP-element group 373: 	393 
    -- CP-element group 373:  members (37) 
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192__exit__
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303__entry__
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Update/cr
      -- 
    crr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1195_call_req_0); -- 
    ccr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1195_call_req_1); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1199_inst_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1208_inst_req_1); -- 
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1218_inst_req_1); -- 
    cr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1228_inst_req_1); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1238_inst_req_1); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1248_inst_req_1); -- 
    cr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1258_inst_req_1); -- 
    cr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1268_inst_req_1); -- 
    cr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1278_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(234) & convTranspose_CP_39_elements(262) & convTranspose_CP_39_elements(296) & convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(364) & convTranspose_CP_39_elements(366) & convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(370) & convTranspose_CP_39_elements(372);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Sample/cra
      -- 
    cra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1195_call_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/call_stmt_1195_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Sample/rr
      -- 
    cca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1195_call_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => type_cast_1199_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Sample/ra
      -- 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	380 
    -- CP-element group 377: 	382 
    -- CP-element group 377: 	384 
    -- CP-element group 377: 	386 
    -- CP-element group 377: 	388 
    -- CP-element group 377: 	390 
    -- CP-element group 377: 	392 
    -- CP-element group 377:  members (27) 
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1199_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Sample/rr
      -- 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    rr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1208_inst_req_0); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1218_inst_req_0); -- 
    rr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1228_inst_req_0); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1238_inst_req_0); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1248_inst_req_0); -- 
    rr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1258_inst_req_0); -- 
    rr_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1268_inst_req_0); -- 
    rr_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1278_inst_req_0); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Sample/ra
      -- 
    ra_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	373 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	414 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1208_Update/ca
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	377 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Sample/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	373 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	411 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1218_Update/ca
      -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Sample/ra
      -- 
    ra_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	373 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	408 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1228_Update/ca
      -- 
    ca_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Sample/ra
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	373 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	405 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1238_Update/ca
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	377 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Sample/ra
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	373 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	402 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1248_Update/ca
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	377 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Sample/ra
      -- 
    ra_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	373 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	399 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1258_Update/ca
      -- 
    ca_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	377 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Sample/ra
      -- 
    ra_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1268_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	373 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	396 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1268_Update/ca
      -- 
    ca_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1268_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	377 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Sample/ra
      -- 
    ra_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1278_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	373 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/type_cast_1278_Update/ca
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Sample/req
      -- 
    ca_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1278_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_0); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Update/req
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_update_start_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Sample/ack
      -- 
    ack_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_1); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Update/ack
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1280_update_completed_
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    -- CP-element group 396:  join  transition  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	391 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Sample/req
      -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_0); -- 
    convTranspose_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(391) & convTranspose_CP_39_elements(395);
      gj_convTranspose_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Sample/ack
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_update_start_
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Update/req
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0, ack => convTranspose_CP_39_elements(397)); -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_1); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1283_Update/ack
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1, ack => convTranspose_CP_39_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	389 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_sample_start_
      -- 
    req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_0); -- 
    convTranspose_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(389) & convTranspose_CP_39_elements(398);
      gj_convTranspose_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Update/req
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_update_start_
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_sample_completed_
      -- 
    ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_1); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1286_update_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	387 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Sample/req
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_sample_start_
      -- 
    req_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_0); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(387) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Update/req
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Sample/ack
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_update_start_
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_sample_completed_
      -- 
    ack_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0, ack => convTranspose_CP_39_elements(403)); -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_1); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Update/ack
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1289_update_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1, ack => convTranspose_CP_39_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	385 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_sample_start_
      -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_0); -- 
    convTranspose_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(385) & convTranspose_CP_39_elements(404);
      gj_convTranspose_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Update/req
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_update_start_
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_sample_completed_
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1292_update_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	383 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_sample_start_
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Sample/req
      -- 
    req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(383) & convTranspose_CP_39_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_update_start_
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Sample/ack
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Update/req
      -- 
    ack_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0, ack => convTranspose_CP_39_elements(409)); -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_1); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1295_Update/ack
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1, ack => convTranspose_CP_39_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	381 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Sample/$entry
      -- 
    req_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_0); -- 
    convTranspose_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(381) & convTranspose_CP_39_elements(410);
      gj_convTranspose_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Update/req
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_update_start_
      -- 
    ack_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0, ack => convTranspose_CP_39_elements(412)); -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_1); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1298_update_completed_
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	379 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_sample_start_
      -- 
    req_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_0); -- 
    convTranspose_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(413);
      gj_convTranspose_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Update/req
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Sample/ack
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_update_start_
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_sample_completed_
      -- 
    ack_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0, ack => convTranspose_CP_39_elements(415)); -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_1); -- 
    -- CP-element group 416:  branch  transition  place  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (13) 
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303__exit__
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305__entry__
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_else_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_if_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_eval_test/branch_req
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_eval_test/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_eval_test/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/if_stmt_1305_dead_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Update/ack
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/R_cmp264505_1306_place
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/WPIPE_ConvTranspose_output_pipe_1301_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1303/$exit
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1, ack => convTranspose_CP_39_elements(416)); -- 
    branch_req_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(416), ack => if_stmt_1305_branch_req_0); -- 
    -- CP-element group 417:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: 	420 
    -- CP-element group 417:  members (18) 
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1311__exit__
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346__entry__
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Update/cr
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Sample/rr
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_update_start_
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/if_stmt_1305_if_link/if_choice_transition
      -- CP-element group 417: 	 branch_block_stmt_32/if_stmt_1305_if_link/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1311_PhiReqMerge
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1311_PhiAck/$entry
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1311_PhiAck/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/merge_stmt_1311_PhiAck/dummy
      -- 
    if_choice_transition_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1305_branch_ack_1, ack => convTranspose_CP_39_elements(417)); -- 
    cr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => type_cast_1332_inst_req_1); -- 
    rr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(417), ack => type_cast_1332_inst_req_0); -- 
    -- CP-element group 418:  transition  place  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	496 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500
      -- CP-element group 418: 	 branch_block_stmt_32/if_stmt_1305_else_link/else_choice_transition
      -- CP-element group 418: 	 branch_block_stmt_32/if_stmt_1305_else_link/$exit
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500_PhiReq/$entry
      -- CP-element group 418: 	 branch_block_stmt_32/forx_xend273_forx_xend500_PhiReq/$exit
      -- 
    else_choice_transition_3080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1305_branch_ack_0, ack => convTranspose_CP_39_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Sample/ra
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_sample_completed_
      -- 
    ra_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_0, ack => convTranspose_CP_39_elements(419)); -- 
    -- CP-element group 420:  transition  place  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	417 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	490 
    -- CP-element group 420:  members (9) 
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346__exit__
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Update/ca
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/type_cast_1332_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1317_to_assign_stmt_1346/$exit
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/$entry
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/$entry
      -- CP-element group 420: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/$entry
      -- 
    ca_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_1, ack => convTranspose_CP_39_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	495 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	466 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Sample/ack
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_sample_complete
      -- 
    ack_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1361_index_offset_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	495 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (11) 
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_offset_calculated
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_root_address_calculated
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_request/req
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_request/$entry
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_base_plus_offset/sum_rename_ack
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_base_plus_offset/sum_rename_req
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_base_plus_offset/$exit
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_base_plus_offset/$entry
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Update/ack
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Update/$exit
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1361_index_offset_ack_1, ack => convTranspose_CP_39_elements(422)); -- 
    req_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => addr_of_1362_final_reg_req_0); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_request/ack
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_request/$exit
      -- 
    ack_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1362_final_reg_ack_0, ack => convTranspose_CP_39_elements(423)); -- 
    -- CP-element group 424:  join  fork  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	495 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (24) 
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_word_addrgen/root_register_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_word_addrgen/root_register_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_word_addrgen/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_word_addrgen/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_plus_offset/sum_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_plus_offset/sum_rename_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_plus_offset/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_plus_offset/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_addr_resize/base_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_addr_resize/base_resize_req
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_addr_resize/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_addr_resize/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_address_resized
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_base_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_complete/ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_complete/$exit
      -- 
    ack_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1362_final_reg_ack_1, ack => convTranspose_CP_39_elements(424)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => ptr_deref_1366_load_0_req_0); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (5) 
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/word_0/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_sample_completed_
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Sample/word_access_start/word_0/ra
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1366_load_0_ack_0, ack => convTranspose_CP_39_elements(425)); -- 
    -- CP-element group 426:  fork  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	495 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426: 	429 
    -- CP-element group 426: 	431 
    -- CP-element group 426: 	433 
    -- CP-element group 426: 	435 
    -- CP-element group 426: 	437 
    -- CP-element group 426: 	439 
    -- CP-element group 426: 	441 
    -- CP-element group 426:  members (33) 
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/ptr_deref_1366_Merge/merge_ack
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/ptr_deref_1366_Merge/merge_req
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/ptr_deref_1366_Merge/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/ptr_deref_1366_Merge/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/word_0/ca
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Sample/$entry
      -- 
    ca_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1366_load_0_ack_1, ack => convTranspose_CP_39_elements(426)); -- 
    rr_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1370_inst_req_0); -- 
    rr_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1380_inst_req_0); -- 
    rr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1390_inst_req_0); -- 
    rr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1400_inst_req_0); -- 
    rr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1410_inst_req_0); -- 
    rr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1420_inst_req_0); -- 
    rr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1430_inst_req_0); -- 
    rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => type_cast_1440_inst_req_0); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Sample/ra
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_sample_completed_
      -- 
    ra_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_0, ack => convTranspose_CP_39_elements(427)); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	495 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	463 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Update/$exit
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Update/ca
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_update_completed_
      -- 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_1, ack => convTranspose_CP_39_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	426 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Sample/ra
      -- 
    ra_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => convTranspose_CP_39_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	495 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	460 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Update/ca
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Update/$exit
      -- 
    ca_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => convTranspose_CP_39_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	426 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Sample/ra
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_sample_completed_
      -- 
    ra_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_0, ack => convTranspose_CP_39_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	495 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	457 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Update/ca
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_update_completed_
      -- 
    ca_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_1, ack => convTranspose_CP_39_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	426 
    -- CP-element group 433: successors 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Sample/ra
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_sample_completed_
      -- 
    ra_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1400_inst_ack_0, ack => convTranspose_CP_39_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	495 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	454 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Update/ca
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_update_completed_
      -- 
    ca_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1400_inst_ack_1, ack => convTranspose_CP_39_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	426 
    -- CP-element group 435: successors 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Sample/ra
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Sample/$exit
      -- 
    ra_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1410_inst_ack_0, ack => convTranspose_CP_39_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	495 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	451 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Update/$exit
      -- 
    ca_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1410_inst_ack_1, ack => convTranspose_CP_39_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	426 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_sample_completed_
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Sample/$exit
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Sample/ra
      -- 
    ra_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1420_inst_ack_0, ack => convTranspose_CP_39_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	495 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	448 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_update_completed_
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Update/ca
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Update/$exit
      -- 
    ca_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1420_inst_ack_1, ack => convTranspose_CP_39_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	426 
    -- CP-element group 439: successors 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Sample/ra
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_sample_completed_
      -- 
    ra_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_0, ack => convTranspose_CP_39_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	495 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	445 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Update/ca
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_update_completed_
      -- 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_1, ack => convTranspose_CP_39_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	426 
    -- CP-element group 441: successors 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Sample/ra
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_sample_completed_
      -- 
    ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1440_inst_ack_0, ack => convTranspose_CP_39_elements(441)); -- 
    -- CP-element group 442:  transition  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	495 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (6) 
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Sample/req
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Update/ca
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_update_completed_
      -- 
    ca_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1440_inst_ack_1, ack => convTranspose_CP_39_elements(442)); -- 
    req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(442), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_0); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Update/req
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Sample/ack
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_update_start_
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_sample_completed_
      -- 
    ack_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0, ack => convTranspose_CP_39_elements(443)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_1); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Update/ack
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1442_update_completed_
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1, ack => convTranspose_CP_39_elements(444)); -- 
    -- CP-element group 445:  join  transition  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	440 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_sample_start_
      -- 
    req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_0); -- 
    convTranspose_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(440) & convTranspose_CP_39_elements(444);
      gj_convTranspose_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Update/req
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Sample/$exit
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_update_start_
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_sample_completed_
      -- 
    ack_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0, ack => convTranspose_CP_39_elements(446)); -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_Update/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1445_update_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	438 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_sample_start_
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Sample/req
      -- CP-element group 448: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Sample/$entry
      -- 
    req_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_0); -- 
    convTranspose_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(438) & convTranspose_CP_39_elements(447);
      gj_convTranspose_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  transition  input  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Update/req
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Sample/ack
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_update_start_
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_sample_completed_
      -- 
    ack_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0, ack => convTranspose_CP_39_elements(449)); -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_1); -- 
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Update/ack
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1448_update_completed_
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1, ack => convTranspose_CP_39_elements(450)); -- 
    -- CP-element group 451:  join  transition  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	436 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Sample/req
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_sample_start_
      -- 
    req_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_0); -- 
    convTranspose_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(436) & convTranspose_CP_39_elements(450);
      gj_convTranspose_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (6) 
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Update/req
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Sample/ack
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_update_start_
      -- CP-element group 452: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_sample_completed_
      -- 
    ack_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0, ack => convTranspose_CP_39_elements(452)); -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_1); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Update/ack
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1451_update_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1, ack => convTranspose_CP_39_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	434 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Sample/req
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_sample_start_
      -- 
    req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(454), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_0); -- 
    convTranspose_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(434) & convTranspose_CP_39_elements(453);
      gj_convTranspose_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  transition  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (6) 
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Sample/ack
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Update/req
      -- 
    ack_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0, ack => convTranspose_CP_39_elements(455)); -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_1); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1454_Update/ack
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1, ack => convTranspose_CP_39_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	432 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Sample/req
      -- 
    req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(457), ack => WPIPE_ConvTranspose_output_pipe_1457_inst_req_0); -- 
    convTranspose_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(432) & convTranspose_CP_39_elements(456);
      gj_convTranspose_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  transition  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (6) 
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_update_start_
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Sample/ack
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Update/req
      -- 
    ack_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0, ack => convTranspose_CP_39_elements(458)); -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1457_inst_req_1); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1457_Update/ack
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1, ack => convTranspose_CP_39_elements(459)); -- 
    -- CP-element group 460:  join  transition  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	430 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Sample/req
      -- 
    req_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(460), ack => WPIPE_ConvTranspose_output_pipe_1460_inst_req_0); -- 
    convTranspose_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(430) & convTranspose_CP_39_elements(459);
      gj_convTranspose_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (6) 
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Sample/ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Update/req
      -- 
    ack_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0, ack => convTranspose_CP_39_elements(461)); -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1460_inst_req_1); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1460_Update/ack
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1, ack => convTranspose_CP_39_elements(462)); -- 
    -- CP-element group 463:  join  transition  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	428 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Sample/req
      -- 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => WPIPE_ConvTranspose_output_pipe_1463_inst_req_0); -- 
    convTranspose_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(428) & convTranspose_CP_39_elements(462);
      gj_convTranspose_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  transition  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (6) 
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_update_start_
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Sample/ack
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Update/$entry
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Update/req
      -- 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1463_inst_req_1); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/WPIPE_ConvTranspose_output_pipe_1463_Update/ack
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1, ack => convTranspose_CP_39_elements(465)); -- 
    -- CP-element group 466:  branch  join  transition  place  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	421 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (10) 
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476__exit__
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477__entry__
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_dead_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_eval_test/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_eval_test/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_eval_test/branch_req
      -- CP-element group 466: 	 branch_block_stmt_32/R_exitcond1_1478_place
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_if_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_32/if_stmt_1477_else_link/$entry
      -- 
    branch_req_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(466), ack => if_stmt_1477_branch_req_0); -- 
    convTranspose_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(421) & convTranspose_CP_39_elements(465);
      gj_convTranspose_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  merge  transition  place  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	496 
    -- CP-element group 467:  members (13) 
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1483__exit__
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500
      -- CP-element group 467: 	 branch_block_stmt_32/if_stmt_1477_if_link/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/if_stmt_1477_if_link/if_choice_transition
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1483_PhiReqMerge
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1483_PhiAck/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1483_PhiAck/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_1483_PhiAck/dummy
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_32/forx_xend500x_xloopexit_forx_xend500_PhiReq/$exit
      -- 
    if_choice_transition_3435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1477_branch_ack_1, ack => convTranspose_CP_39_elements(467)); -- 
    -- CP-element group 468:  fork  transition  place  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	491 
    -- CP-element group 468: 	492 
    -- CP-element group 468:  members (12) 
      -- CP-element group 468: 	 branch_block_stmt_32/if_stmt_1477_else_link/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/if_stmt_1477_else_link/else_choice_transition
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Sample/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Sample/rr
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1477_branch_ack_0, ack => convTranspose_CP_39_elements(468)); -- 
    rr_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => type_cast_1355_inst_req_0); -- 
    cr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => type_cast_1355_inst_req_1); -- 
    -- CP-element group 469:  merge  branch  transition  place  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	165 
    -- CP-element group 469: 	120 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	121 
    -- CP-element group 469: 	122 
    -- CP-element group 469:  members (17) 
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424__exit__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430__entry__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430__exit__
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431__entry__
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_430/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_dead_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_eval_test/branch_req
      -- CP-element group 469: 	 branch_block_stmt_32/R_cmp194509_432_place
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_if_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/if_stmt_431_else_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiReqMerge
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/dummy
      -- 
    branch_req_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => if_stmt_431_branch_req_0); -- 
    convTranspose_CP_39_elements(469) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 470:  transition  output  delay-element  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	124 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	474 
    -- CP-element group 470:  members (5) 
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_473_konst_delay_trans
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- 
    phi_stmt_469_req_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(470), ack => phi_stmt_469_req_0); -- 
    -- Element group convTranspose_CP_39_elements(470) is a control-delay.
    cp_element_470_delay: control_delay_element  generic map(name => " 470_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(470), clk => clk, reset =>reset);
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	166 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (2) 
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/ra
      -- 
    ra_3507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_0, ack => convTranspose_CP_39_elements(471)); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	166 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/ca
      -- 
    ca_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_1, ack => convTranspose_CP_39_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (6) 
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- 
    phi_stmt_469_req_3513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(473), ack => phi_stmt_469_req_1); -- 
    convTranspose_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(471) & convTranspose_CP_39_elements(472);
      gj_convTranspose_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  merge  transition  place  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	470 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (2) 
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_468_PhiReqMerge
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(474) <= OrReduce(convTranspose_CP_39_elements(470) & convTranspose_CP_39_elements(473));
    -- CP-element group 475:  fork  transition  place  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	163 
    -- CP-element group 475: 	156 
    -- CP-element group 475: 	160 
    -- CP-element group 475: 	152 
    -- CP-element group 475: 	125 
    -- CP-element group 475: 	126 
    -- CP-element group 475: 	128 
    -- CP-element group 475: 	129 
    -- CP-element group 475: 	132 
    -- CP-element group 475: 	136 
    -- CP-element group 475: 	140 
    -- CP-element group 475: 	144 
    -- CP-element group 475: 	148 
    -- CP-element group 475:  members (56) 
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468__exit__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__entry__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resized_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scaled_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_computed_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_update_start
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/rr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/phi_stmt_469_ack
      -- 
    phi_stmt_469_ack_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_469_ack_0, ack => convTranspose_CP_39_elements(475)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_538_inst_req_1); -- 
    cr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => ptr_deref_618_store_0_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_610_inst_req_1); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_574_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_556_inst_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_592_inst_req_1); -- 
    req_981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_481_index_offset_req_0); -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_481_index_offset_req_1); -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => addr_of_482_final_reg_req_1); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_0); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_489_inst_req_1); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_502_inst_req_1); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_520_inst_req_1); -- 
    -- CP-element group 476:  transition  output  delay-element  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	168 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	480 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_682_konst_delay_trans
      -- CP-element group 476: 	 branch_block_stmt_32/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(476), ack => phi_stmt_676_req_1); -- 
    -- Element group convTranspose_CP_39_elements(476) is a control-delay.
    cp_element_476_delay: control_delay_element  generic map(name => " 476_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(476), clk => clk, reset =>reset);
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	210 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (2) 
      -- CP-element group 477: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$exit
      -- CP-element group 477: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/ra
      -- 
    ra_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => convTranspose_CP_39_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	210 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/ca
      -- 
    ca_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => convTranspose_CP_39_elements(478)); -- 
    -- CP-element group 479:  join  transition  output  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: 	478 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (6) 
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(479), ack => phi_stmt_676_req_0); -- 
    convTranspose_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(477) & convTranspose_CP_39_elements(478);
      gj_convTranspose_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  merge  transition  place  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	476 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (2) 
      -- CP-element group 480: 	 branch_block_stmt_32/merge_stmt_675_PhiReqMerge
      -- CP-element group 480: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(480) <= OrReduce(convTranspose_CP_39_elements(476) & convTranspose_CP_39_elements(479));
    -- CP-element group 481:  fork  transition  place  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	169 
    -- CP-element group 481: 	170 
    -- CP-element group 481: 	172 
    -- CP-element group 481: 	173 
    -- CP-element group 481: 	176 
    -- CP-element group 481: 	180 
    -- CP-element group 481: 	184 
    -- CP-element group 481: 	188 
    -- CP-element group 481: 	192 
    -- CP-element group 481: 	196 
    -- CP-element group 481: 	200 
    -- CP-element group 481: 	204 
    -- CP-element group 481: 	207 
    -- CP-element group 481:  members (56) 
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675__exit__
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__entry__
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resized_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_update_start
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_ack
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_ack
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_req
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_computed_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scaled_1
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/cr
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/phi_stmt_676_ack
      -- 
    phi_stmt_676_ack_3572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_676_ack_0, ack => convTranspose_CP_39_elements(481)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_727_inst_req_1); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_709_inst_req_1); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => addr_of_689_final_reg_req_1); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_0); -- 
    req_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => array_obj_ref_688_index_offset_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_696_inst_req_1); -- 
    req_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => array_obj_ref_688_index_offset_req_0); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_745_inst_req_1); -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_763_inst_req_1); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_781_inst_req_1); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_799_inst_req_1); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => type_cast_817_inst_req_1); -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => ptr_deref_825_store_0_req_1); -- 
    -- CP-element group 482:  merge  fork  transition  place  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	209 
    -- CP-element group 482: 	122 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	211 
    -- CP-element group 482: 	212 
    -- CP-element group 482: 	213 
    -- CP-element group 482: 	214 
    -- CP-element group 482: 	215 
    -- CP-element group 482: 	216 
    -- CP-element group 482:  members (25) 
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847__exit__
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__entry__
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiReqMerge
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/dummy
      -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_850_inst_req_0); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_850_inst_req_1); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_854_inst_req_0); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_854_inst_req_1); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_858_inst_req_0); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => type_cast_858_inst_req_1); -- 
    convTranspose_CP_39_elements(482) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 483:  transition  output  delay-element  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	221 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	487 
    -- CP-element group 483:  members (5) 
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_926_konst_delay_trans
      -- CP-element group 483: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(483), ack => phi_stmt_920_req_1); -- 
    -- Element group convTranspose_CP_39_elements(483) is a control-delay.
    cp_element_483_delay: control_delay_element  generic map(name => " 483_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(483), clk => clk, reset =>reset);
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	230 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	486 
    -- CP-element group 484:  members (2) 
      -- CP-element group 484: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/ra
      -- 
    ra_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => convTranspose_CP_39_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	230 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (2) 
      -- CP-element group 485: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/ca
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => convTranspose_CP_39_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	484 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (6) 
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(486), ack => phi_stmt_920_req_0); -- 
    convTranspose_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(484) & convTranspose_CP_39_elements(485);
      gj_convTranspose_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  merge  transition  place  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	483 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (2) 
      -- CP-element group 487: 	 branch_block_stmt_32/merge_stmt_919_PhiReqMerge
      -- CP-element group 487: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(487) <= OrReduce(convTranspose_CP_39_elements(483) & convTranspose_CP_39_elements(486));
    -- CP-element group 488:  fork  transition  place  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	222 
    -- CP-element group 488: 	223 
    -- CP-element group 488: 	225 
    -- CP-element group 488: 	227 
    -- CP-element group 488:  members (29) 
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919__exit__
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__entry__
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_start_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resized_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scaled_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_computed_1
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_ack
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_ack
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_update_start
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/req
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_start_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/cr
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/phi_stmt_920_ack
      -- 
    phi_stmt_920_ack_3649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_920_ack_0, ack => convTranspose_CP_39_elements(488)); -- 
    req_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => array_obj_ref_932_index_offset_req_0); -- 
    req_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => array_obj_ref_932_index_offset_req_1); -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => addr_of_933_final_reg_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => ptr_deref_936_store_0_req_1); -- 
    -- CP-element group 489:  merge  fork  transition  place  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	219 
    -- CP-element group 489: 	229 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	231 
    -- CP-element group 489: 	232 
    -- CP-element group 489: 	234 
    -- CP-element group 489: 	235 
    -- CP-element group 489: 	263 
    -- CP-element group 489: 	281 
    -- CP-element group 489: 	282 
    -- CP-element group 489: 	286 
    -- CP-element group 489: 	287 
    -- CP-element group 489: 	297 
    -- CP-element group 489: 	315 
    -- CP-element group 489: 	316 
    -- CP-element group 489: 	320 
    -- CP-element group 489: 	321 
    -- CP-element group 489: 	331 
    -- CP-element group 489: 	349 
    -- CP-element group 489: 	350 
    -- CP-element group 489: 	354 
    -- CP-element group 489: 	355 
    -- CP-element group 489: 	365 
    -- CP-element group 489: 	367 
    -- CP-element group 489: 	369 
    -- CP-element group 489: 	371 
    -- CP-element group 489:  members (76) 
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959__exit__
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192__entry__
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/crr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/ccr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_update_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/rr
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiReqMerge
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$entry
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$exit
      -- CP-element group 489: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/dummy
      -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1048_inst_req_0); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => WPIPE_Block1_start_1013_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1048_inst_req_1); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => WPIPE_Block2_start_1069_inst_req_0); -- 
    cr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1055_inst_req_1); -- 
    rr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1055_inst_req_0); -- 
    crr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => call_stmt_962_call_req_0); -- 
    ccr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => call_stmt_962_call_req_1); -- 
    cr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_967_inst_req_1); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => WPIPE_Block0_start_969_inst_req_0); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1104_inst_req_0); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1104_inst_req_1); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1111_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1111_inst_req_1); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => WPIPE_Block3_start_1125_inst_req_0); -- 
    rr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1160_inst_req_0); -- 
    cr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1160_inst_req_1); -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1167_inst_req_0); -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => type_cast_1167_inst_req_1); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => RPIPE_Block0_done_1182_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => RPIPE_Block1_done_1185_inst_req_0); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => RPIPE_Block2_done_1188_inst_req_0); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(489), ack => RPIPE_Block3_done_1191_inst_req_0); -- 
    convTranspose_CP_39_elements(489) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 490:  transition  output  delay-element  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	420 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	494 
    -- CP-element group 490:  members (5) 
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/$exit
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1353_konst_delay_trans
      -- CP-element group 490: 	 branch_block_stmt_32/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_req
      -- 
    phi_stmt_1349_req_3695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1349_req_3695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(490), ack => phi_stmt_1349_req_0); -- 
    -- Element group convTranspose_CP_39_elements(490) is a control-delay.
    cp_element_490_delay: control_delay_element  generic map(name => " 490_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(420), ack => convTranspose_CP_39_elements(490), clk => clk, reset =>reset);
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	468 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (2) 
      -- CP-element group 491: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Sample/ra
      -- 
    ra_3715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_0, ack => convTranspose_CP_39_elements(491)); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	468 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (2) 
      -- CP-element group 492: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/Update/ca
      -- 
    ca_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_1, ack => convTranspose_CP_39_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (6) 
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_sources/type_cast_1355/SplitProtocol/$exit
      -- CP-element group 493: 	 branch_block_stmt_32/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1349/phi_stmt_1349_req
      -- 
    phi_stmt_1349_req_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1349_req_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(493), ack => phi_stmt_1349_req_1); -- 
    convTranspose_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(491) & convTranspose_CP_39_elements(492);
      gj_convTranspose_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  merge  transition  place  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	490 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (2) 
      -- CP-element group 494: 	 branch_block_stmt_32/merge_stmt_1348_PhiReqMerge
      -- CP-element group 494: 	 branch_block_stmt_32/merge_stmt_1348_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(494) <= OrReduce(convTranspose_CP_39_elements(490) & convTranspose_CP_39_elements(493));
    -- CP-element group 495:  fork  transition  place  input  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	421 
    -- CP-element group 495: 	422 
    -- CP-element group 495: 	424 
    -- CP-element group 495: 	426 
    -- CP-element group 495: 	428 
    -- CP-element group 495: 	430 
    -- CP-element group 495: 	432 
    -- CP-element group 495: 	434 
    -- CP-element group 495: 	436 
    -- CP-element group 495: 	438 
    -- CP-element group 495: 	440 
    -- CP-element group 495: 	442 
    -- CP-element group 495:  members (53) 
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_resize_1/index_resize_req
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1348__exit__
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476__entry__
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_resized_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_resize_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_resize_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_scaled_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1400_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1370_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/word_0/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_complete/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/word_0/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/addr_of_1362_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_computed_1
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1390_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1440_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1410_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Update/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/word_access_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Sample/req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/ptr_deref_1366_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_final_index_sum_regn_update_start
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_scale_1/scale_rename_ack
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1430_update_start_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_scale_1/scale_rename_req
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_scale_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1380_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_scale_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/array_obj_ref_1361_index_resize_1/index_resize_ack
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1363_to_assign_stmt_1476/type_cast_1420_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1348_PhiAck/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/merge_stmt_1348_PhiAck/phi_stmt_1349_ack
      -- 
    phi_stmt_1349_ack_3726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1349_ack_0, ack => convTranspose_CP_39_elements(495)); -- 
    cr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1400_inst_req_1); -- 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1370_inst_req_1); -- 
    cr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1410_inst_req_1); -- 
    cr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1390_inst_req_1); -- 
    cr_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => ptr_deref_1366_load_0_req_1); -- 
    req_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => addr_of_1362_final_reg_req_1); -- 
    cr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1440_inst_req_1); -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => array_obj_ref_1361_index_offset_req_1); -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1430_inst_req_1); -- 
    req_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => array_obj_ref_1361_index_offset_req_0); -- 
    cr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1380_inst_req_1); -- 
    cr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(495), ack => type_cast_1420_inst_req_1); -- 
    -- CP-element group 496:  merge  transition  place  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	418 
    -- CP-element group 496: 	467 
    -- CP-element group 496: successors 
    -- CP-element group 496:  members (16) 
      -- CP-element group 496: 	 $exit
      -- CP-element group 496: 	 branch_block_stmt_32/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1485__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/return__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1487__exit__
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1485_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1485_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1485_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1485_PhiAck/dummy
      -- CP-element group 496: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1487_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1487_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1487_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_32/merge_stmt_1487_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(496) <= OrReduce(convTranspose_CP_39_elements(418) & convTranspose_CP_39_elements(467));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar525_931_resized : std_logic_vector(13 downto 0);
    signal R_indvar525_931_scaled : std_logic_vector(13 downto 0);
    signal R_indvar539_687_resized : std_logic_vector(10 downto 0);
    signal R_indvar539_687_scaled : std_logic_vector(10 downto 0);
    signal R_indvar555_480_resized : std_logic_vector(13 downto 0);
    signal R_indvar555_480_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1360_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1360_scaled : std_logic_vector(13 downto 0);
    signal add108_333 : std_logic_vector(15 downto 0);
    signal add117_358 : std_logic_vector(15 downto 0);
    signal add126_383 : std_logic_vector(15 downto 0);
    signal add12_82 : std_logic_vector(15 downto 0);
    signal add135_408 : std_logic_vector(15 downto 0);
    signal add150_508 : std_logic_vector(63 downto 0);
    signal add156_526 : std_logic_vector(63 downto 0);
    signal add162_544 : std_logic_vector(63 downto 0);
    signal add168_562 : std_logic_vector(63 downto 0);
    signal add174_580 : std_logic_vector(63 downto 0);
    signal add180_598 : std_logic_vector(63 downto 0);
    signal add186_616 : std_logic_vector(63 downto 0);
    signal add206_715 : std_logic_vector(63 downto 0);
    signal add212_733 : std_logic_vector(63 downto 0);
    signal add218_751 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(15 downto 0);
    signal add224_769 : std_logic_vector(63 downto 0);
    signal add230_787 : std_logic_vector(63 downto 0);
    signal add236_805 : std_logic_vector(63 downto 0);
    signal add242_823 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(15 downto 0);
    signal add39_157 : std_logic_vector(15 downto 0);
    signal add48_182 : std_logic_vector(15 downto 0);
    signal add57_207 : std_logic_vector(15 downto 0);
    signal add74_247 : std_logic_vector(31 downto 0);
    signal add79_252 : std_logic_vector(31 downto 0);
    signal add99_308 : std_logic_vector(15 downto 0);
    signal add_57 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1361_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1361_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1361_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1361_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1361_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1361_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_688_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_932_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_690 : std_logic_vector(31 downto 0);
    signal arrayidx269_934 : std_logic_vector(31 downto 0);
    signal arrayidx432_1363 : std_logic_vector(31 downto 0);
    signal arrayidx_483 : std_logic_vector(31 downto 0);
    signal call101_311 : std_logic_vector(7 downto 0);
    signal call106_324 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_336 : std_logic_vector(7 downto 0);
    signal call115_349 : std_logic_vector(7 downto 0);
    signal call119_361 : std_logic_vector(7 downto 0);
    signal call124_374 : std_logic_vector(7 downto 0);
    signal call128_386 : std_logic_vector(7 downto 0);
    signal call133_399 : std_logic_vector(7 downto 0);
    signal call143_486 : std_logic_vector(7 downto 0);
    signal call147_499 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_517 : std_logic_vector(7 downto 0);
    signal call159_535 : std_logic_vector(7 downto 0);
    signal call165_553 : std_logic_vector(7 downto 0);
    signal call171_571 : std_logic_vector(7 downto 0);
    signal call177_589 : std_logic_vector(7 downto 0);
    signal call183_607 : std_logic_vector(7 downto 0);
    signal call199_693 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_706 : std_logic_vector(7 downto 0);
    signal call209_724 : std_logic_vector(7 downto 0);
    signal call215_742 : std_logic_vector(7 downto 0);
    signal call221_760 : std_logic_vector(7 downto 0);
    signal call227_778 : std_logic_vector(7 downto 0);
    signal call233_796 : std_logic_vector(7 downto 0);
    signal call239_814 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_962 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call346_1183 : std_logic_vector(15 downto 0);
    signal call348_1186 : std_logic_vector(15 downto 0);
    signal call350_1189 : std_logic_vector(15 downto 0);
    signal call352_1192 : std_logic_vector(15 downto 0);
    signal call354_1195 : std_logic_vector(63 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call92_286 : std_logic_vector(7 downto 0);
    signal call97_299 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194509_430 : std_logic_vector(0 downto 0);
    signal cmp264505_875 : std_logic_vector(0 downto 0);
    signal cmp513_415 : std_logic_vector(0 downto 0);
    signal conv104_315 : std_logic_vector(15 downto 0);
    signal conv107_328 : std_logic_vector(15 downto 0);
    signal conv113_340 : std_logic_vector(15 downto 0);
    signal conv116_353 : std_logic_vector(15 downto 0);
    signal conv11_77 : std_logic_vector(15 downto 0);
    signal conv122_365 : std_logic_vector(15 downto 0);
    signal conv125_378 : std_logic_vector(15 downto 0);
    signal conv131_390 : std_logic_vector(15 downto 0);
    signal conv134_403 : std_logic_vector(15 downto 0);
    signal conv144_490 : std_logic_vector(63 downto 0);
    signal conv149_503 : std_logic_vector(63 downto 0);
    signal conv155_521 : std_logic_vector(63 downto 0);
    signal conv161_539 : std_logic_vector(63 downto 0);
    signal conv167_557 : std_logic_vector(63 downto 0);
    signal conv173_575 : std_logic_vector(63 downto 0);
    signal conv179_593 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(15 downto 0);
    signal conv185_611 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(15 downto 0);
    signal conv200_697 : std_logic_vector(63 downto 0);
    signal conv205_710 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(15 downto 0);
    signal conv211_728 : std_logic_vector(63 downto 0);
    signal conv217_746 : std_logic_vector(63 downto 0);
    signal conv223_764 : std_logic_vector(63 downto 0);
    signal conv229_782 : std_logic_vector(63 downto 0);
    signal conv235_800 : std_logic_vector(63 downto 0);
    signal conv241_818 : std_logic_vector(63 downto 0);
    signal conv253_851 : std_logic_vector(31 downto 0);
    signal conv255_855 : std_logic_vector(31 downto 0);
    signal conv258_859 : std_logic_vector(31 downto 0);
    signal conv26_114 : std_logic_vector(15 downto 0);
    signal conv276_968 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(15 downto 0);
    signal conv305_1049 : std_logic_vector(15 downto 0);
    signal conv307_1056 : std_logic_vector(15 downto 0);
    signal conv322_1105 : std_logic_vector(15 downto 0);
    signal conv324_1112 : std_logic_vector(15 downto 0);
    signal conv339_1161 : std_logic_vector(15 downto 0);
    signal conv341_1168 : std_logic_vector(15 downto 0);
    signal conv355_1200 : std_logic_vector(63 downto 0);
    signal conv35_139 : std_logic_vector(15 downto 0);
    signal conv361_1209 : std_logic_vector(7 downto 0);
    signal conv367_1219 : std_logic_vector(7 downto 0);
    signal conv373_1229 : std_logic_vector(7 downto 0);
    signal conv379_1239 : std_logic_vector(7 downto 0);
    signal conv385_1249 : std_logic_vector(7 downto 0);
    signal conv38_152 : std_logic_vector(15 downto 0);
    signal conv391_1259 : std_logic_vector(7 downto 0);
    signal conv397_1269 : std_logic_vector(7 downto 0);
    signal conv3_52 : std_logic_vector(15 downto 0);
    signal conv403_1279 : std_logic_vector(7 downto 0);
    signal conv437_1371 : std_logic_vector(7 downto 0);
    signal conv443_1381 : std_logic_vector(7 downto 0);
    signal conv449_1391 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(15 downto 0);
    signal conv455_1401 : std_logic_vector(7 downto 0);
    signal conv461_1411 : std_logic_vector(7 downto 0);
    signal conv467_1421 : std_logic_vector(7 downto 0);
    signal conv473_1431 : std_logic_vector(7 downto 0);
    signal conv479_1441 : std_logic_vector(7 downto 0);
    signal conv47_177 : std_logic_vector(15 downto 0);
    signal conv53_189 : std_logic_vector(15 downto 0);
    signal conv56_202 : std_logic_vector(15 downto 0);
    signal conv61_211 : std_logic_vector(31 downto 0);
    signal conv63_215 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv82_256 : std_logic_vector(31 downto 0);
    signal conv84_260 : std_logic_vector(31 downto 0);
    signal conv87_264 : std_logic_vector(31 downto 0);
    signal conv8_64 : std_logic_vector(15 downto 0);
    signal conv90_268 : std_logic_vector(31 downto 0);
    signal conv95_290 : std_logic_vector(15 downto 0);
    signal conv98_303 : std_logic_vector(15 downto 0);
    signal exitcond1_1476 : std_logic_vector(0 downto 0);
    signal exitcond2_838 : std_logic_vector(0 downto 0);
    signal exitcond3_631 : std_logic_vector(0 downto 0);
    signal exitcond_950 : std_logic_vector(0 downto 0);
    signal iNsTr_14_241 : std_logic_vector(31 downto 0);
    signal iNsTr_194_1333 : std_logic_vector(63 downto 0);
    signal iNsTr_26_453 : std_logic_vector(63 downto 0);
    signal iNsTr_39_660 : std_logic_vector(63 downto 0);
    signal iNsTr_53_904 : std_logic_vector(63 downto 0);
    signal indvar525_920 : std_logic_vector(63 downto 0);
    signal indvar539_676 : std_logic_vector(63 downto 0);
    signal indvar555_469 : std_logic_vector(63 downto 0);
    signal indvar_1349 : std_logic_vector(63 downto 0);
    signal indvarx_xnext526_945 : std_logic_vector(63 downto 0);
    signal indvarx_xnext540_833 : std_logic_vector(63 downto 0);
    signal indvarx_xnext556_626 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1471 : std_logic_vector(63 downto 0);
    signal mul256_864 : std_logic_vector(31 downto 0);
    signal mul259_869 : std_logic_vector(31 downto 0);
    signal mul66_229 : std_logic_vector(31 downto 0);
    signal mul85_273 : std_logic_vector(31 downto 0);
    signal mul88_278 : std_logic_vector(31 downto 0);
    signal mul91_283 : std_logic_vector(31 downto 0);
    signal mul_224 : std_logic_vector(31 downto 0);
    signal ptr_deref_1366_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1366_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1366_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1366_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1366_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_618_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_618_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_825_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_825_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_825_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_825_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_936_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_936_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_936_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_936_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_321 : std_logic_vector(15 downto 0);
    signal shl114_346 : std_logic_vector(15 downto 0);
    signal shl123_371 : std_logic_vector(15 downto 0);
    signal shl132_396 : std_logic_vector(15 downto 0);
    signal shl146_496 : std_logic_vector(63 downto 0);
    signal shl152_514 : std_logic_vector(63 downto 0);
    signal shl158_532 : std_logic_vector(63 downto 0);
    signal shl164_550 : std_logic_vector(63 downto 0);
    signal shl170_568 : std_logic_vector(63 downto 0);
    signal shl176_586 : std_logic_vector(63 downto 0);
    signal shl182_604 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(15 downto 0);
    signal shl202_703 : std_logic_vector(63 downto 0);
    signal shl208_721 : std_logic_vector(63 downto 0);
    signal shl214_739 : std_logic_vector(63 downto 0);
    signal shl220_757 : std_logic_vector(63 downto 0);
    signal shl226_775 : std_logic_vector(63 downto 0);
    signal shl232_793 : std_logic_vector(63 downto 0);
    signal shl238_811 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(15 downto 0);
    signal shl36_145 : std_logic_vector(15 downto 0);
    signal shl45_170 : std_logic_vector(15 downto 0);
    signal shl54_195 : std_logic_vector(15 downto 0);
    signal shl96_296 : std_logic_vector(15 downto 0);
    signal shl9_70 : std_logic_vector(15 downto 0);
    signal shl_45 : std_logic_vector(15 downto 0);
    signal shr304_1045 : std_logic_vector(31 downto 0);
    signal shr321_1101 : std_logic_vector(31 downto 0);
    signal shr338_1157 : std_logic_vector(31 downto 0);
    signal shr364_1215 : std_logic_vector(63 downto 0);
    signal shr370_1225 : std_logic_vector(63 downto 0);
    signal shr376_1235 : std_logic_vector(63 downto 0);
    signal shr382_1245 : std_logic_vector(63 downto 0);
    signal shr388_1255 : std_logic_vector(63 downto 0);
    signal shr394_1265 : std_logic_vector(63 downto 0);
    signal shr400_1275 : std_logic_vector(63 downto 0);
    signal shr440_1377 : std_logic_vector(63 downto 0);
    signal shr446_1387 : std_logic_vector(63 downto 0);
    signal shr452_1397 : std_logic_vector(63 downto 0);
    signal shr458_1407 : std_logic_vector(63 downto 0);
    signal shr464_1417 : std_logic_vector(63 downto 0);
    signal shr470_1427 : std_logic_vector(63 downto 0);
    signal shr476_1437 : std_logic_vector(63 downto 0);
    signal shr_235 : std_logic_vector(31 downto 0);
    signal sub_1205 : std_logic_vector(63 downto 0);
    signal tmp433_1367 : std_logic_vector(63 downto 0);
    signal tmp520_1317 : std_logic_vector(31 downto 0);
    signal tmp520x_xop_1329 : std_logic_vector(31 downto 0);
    signal tmp521_1323 : std_logic_vector(0 downto 0);
    signal tmp524_1346 : std_logic_vector(63 downto 0);
    signal tmp532_888 : std_logic_vector(31 downto 0);
    signal tmp532x_xop_900 : std_logic_vector(31 downto 0);
    signal tmp533_894 : std_logic_vector(0 downto 0);
    signal tmp537_917 : std_logic_vector(63 downto 0);
    signal tmp548_644 : std_logic_vector(31 downto 0);
    signal tmp548x_xop_656 : std_logic_vector(31 downto 0);
    signal tmp549_650 : std_logic_vector(0 downto 0);
    signal tmp553_673 : std_logic_vector(63 downto 0);
    signal tmp562x_xop_449 : std_logic_vector(31 downto 0);
    signal tmp563_443 : std_logic_vector(0 downto 0);
    signal tmp567_466 : std_logic_vector(63 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1043_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1155_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1198_wire : std_logic_vector(63 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1223_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1253_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1263_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1273_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1315_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1321_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1327_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1337_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1355_wire : std_logic_vector(63 downto 0);
    signal type_cast_1375_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1385_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1395_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1405_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1415_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1425_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1435_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1469_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_294_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_319_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_475_wire : std_logic_vector(63 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_602_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_671_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_679_wire : std_logic_vector(63 downto 0);
    signal type_cast_682_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_923_wire : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_966_wire : std_logic_vector(63 downto 0);
    signal type_cast_998_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop569_910 : std_logic_vector(63 downto 0);
    signal xx_xop570_666 : std_logic_vector(63 downto 0);
    signal xx_xop571_459 : std_logic_vector(63 downto 0);
    signal xx_xop_1339 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1361_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1361_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1361_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1361_resized_base_address <= "00000000000000";
    array_obj_ref_481_constant_part_of_offset <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_481_resized_base_address <= "00000000000000";
    array_obj_ref_688_constant_part_of_offset <= "00000100010";
    array_obj_ref_688_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_688_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_688_resized_base_address <= "00000000000";
    array_obj_ref_932_constant_part_of_offset <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_932_resized_base_address <= "00000000000000";
    ptr_deref_1366_word_offset_0 <= "00000000000000";
    ptr_deref_618_word_offset_0 <= "00000000000000";
    ptr_deref_825_word_offset_0 <= "00000000000";
    ptr_deref_936_word_offset_0 <= "00000000000000";
    type_cast_1002_wire_constant <= "0000000000000000";
    type_cast_1043_wire_constant <= "00000000000000000000000000010010";
    type_cast_1099_wire_constant <= "00000000000000000000000000010001";
    type_cast_1155_wire_constant <= "00000000000000000000000000010000";
    type_cast_118_wire_constant <= "0000000000001000";
    type_cast_1213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1223_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1233_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1243_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1253_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1263_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1273_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1315_wire_constant <= "00000000000000000000000000000010";
    type_cast_1321_wire_constant <= "00000000000000000000000000000001";
    type_cast_1327_wire_constant <= "11111111111111111111111111111111";
    type_cast_1337_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1344_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1375_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1385_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1405_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1415_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1425_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1435_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_143_wire_constant <= "0000000000001000";
    type_cast_1469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_168_wire_constant <= "0000000000001000";
    type_cast_193_wire_constant <= "0000000000001000";
    type_cast_233_wire_constant <= "00000000000000000000000000000010";
    type_cast_239_wire_constant <= "00000000000000000000000000000001";
    type_cast_245_wire_constant <= "01111111111111111111111111111110";
    type_cast_294_wire_constant <= "0000000000001000";
    type_cast_319_wire_constant <= "0000000000001000";
    type_cast_344_wire_constant <= "0000000000001000";
    type_cast_369_wire_constant <= "0000000000001000";
    type_cast_394_wire_constant <= "0000000000001000";
    type_cast_412_wire_constant <= "00000000000000000000000000000011";
    type_cast_428_wire_constant <= "00000000000000000000000000000011";
    type_cast_43_wire_constant <= "0000000000001000";
    type_cast_441_wire_constant <= "00000000000000000000000000000001";
    type_cast_447_wire_constant <= "11111111111111111111111111111111";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_494_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_584_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_602_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_642_wire_constant <= "00000000000000000000000000000010";
    type_cast_648_wire_constant <= "00000000000000000000000000000001";
    type_cast_654_wire_constant <= "11111111111111111111111111111111";
    type_cast_664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_671_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_682_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_68_wire_constant <= "0000000000001000";
    type_cast_701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_737_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_791_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_831_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_873_wire_constant <= "00000000000000000000000000000011";
    type_cast_886_wire_constant <= "00000000000000000000000000000010";
    type_cast_892_wire_constant <= "00000000000000000000000000000001";
    type_cast_898_wire_constant <= "11111111111111111111111111111111";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_915_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_938_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_93_wire_constant <= "0000000000001000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_998_wire_constant <= "0000000000000000";
    phi_stmt_1349: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1353_wire_constant & type_cast_1355_wire;
      req <= phi_stmt_1349_req_0 & phi_stmt_1349_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1349",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1349_ack_0,
          idata => idata,
          odata => indvar_1349,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1349
    phi_stmt_469: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_473_wire_constant & type_cast_475_wire;
      req <= phi_stmt_469_req_0 & phi_stmt_469_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_469",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_469_ack_0,
          idata => idata,
          odata => indvar555_469,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_469
    phi_stmt_676: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_679_wire & type_cast_682_wire_constant;
      req <= phi_stmt_676_req_0 & phi_stmt_676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_676",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_676_ack_0,
          idata => idata,
          odata => indvar539_676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_676
    phi_stmt_920: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_923_wire & type_cast_926_wire_constant;
      req <= phi_stmt_920_req_0 & phi_stmt_920_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_920",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_920_ack_0,
          idata => idata,
          odata => indvar525_920,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_920
    -- flow-through select operator MUX_1345_inst
    tmp524_1346 <= xx_xop_1339 when (tmp521_1323(0) /=  '0') else type_cast_1344_wire_constant;
    -- flow-through select operator MUX_465_inst
    tmp567_466 <= xx_xop571_459 when (tmp563_443(0) /=  '0') else type_cast_464_wire_constant;
    -- flow-through select operator MUX_672_inst
    tmp553_673 <= xx_xop570_666 when (tmp549_650(0) /=  '0') else type_cast_671_wire_constant;
    -- flow-through select operator MUX_916_inst
    tmp537_917 <= xx_xop569_910 when (tmp533_894(0) /=  '0') else type_cast_915_wire_constant;
    addr_of_1362_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1362_final_reg_req_0;
      addr_of_1362_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1362_final_reg_req_1;
      addr_of_1362_final_reg_ack_1<= rack(0);
      addr_of_1362_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1362_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1361_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx432_1363,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_482_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_482_final_reg_req_0;
      addr_of_482_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_482_final_reg_req_1;
      addr_of_482_final_reg_ack_1<= rack(0);
      addr_of_482_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_482_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_481_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_689_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_689_final_reg_req_0;
      addr_of_689_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_689_final_reg_req_1;
      addr_of_689_final_reg_ack_1<= rack(0);
      addr_of_689_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_689_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_688_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_933_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_933_final_reg_req_0;
      addr_of_933_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_933_final_reg_req_1;
      addr_of_933_final_reg_ack_1<= rack(0);
      addr_of_933_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_933_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_932_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1048_inst_req_0;
      type_cast_1048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1048_inst_req_1;
      type_cast_1048_inst_ack_1<= rack(0);
      type_cast_1048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1160_inst_req_0;
      type_cast_1160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1160_inst_req_1;
      type_cast_1160_inst_ack_1<= rack(0);
      type_cast_1160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1199_inst_req_0;
      type_cast_1199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1199_inst_req_1;
      type_cast_1199_inst_ack_1<= rack(0);
      type_cast_1199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1198_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1208_inst_req_0;
      type_cast_1208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1208_inst_req_1;
      type_cast_1208_inst_ack_1<= rack(0);
      type_cast_1208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1218_inst_req_0;
      type_cast_1218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1218_inst_req_1;
      type_cast_1218_inst_ack_1<= rack(0);
      type_cast_1218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1228_inst_req_0;
      type_cast_1228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1228_inst_req_1;
      type_cast_1228_inst_ack_1<= rack(0);
      type_cast_1228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1248_inst_req_0;
      type_cast_1248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1248_inst_req_1;
      type_cast_1248_inst_ack_1<= rack(0);
      type_cast_1248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr382_1245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_1249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1258_inst_req_0;
      type_cast_1258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1258_inst_req_1;
      type_cast_1258_inst_ack_1<= rack(0);
      type_cast_1258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr388_1255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1268_inst_req_0;
      type_cast_1268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1268_inst_req_1;
      type_cast_1268_inst_ack_1<= rack(0);
      type_cast_1268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr394_1265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_1269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1278_inst_req_0;
      type_cast_1278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1278_inst_req_1;
      type_cast_1278_inst_ack_1<= rack(0);
      type_cast_1278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr400_1275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv403_1279,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1332_inst_req_0;
      type_cast_1332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1332_inst_req_1;
      type_cast_1332_inst_ack_1<= rack(0);
      type_cast_1332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp520x_xop_1329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_194_1333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1355_inst_req_0;
      type_cast_1355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1355_inst_req_1;
      type_cast_1355_inst_ack_1<= rack(0);
      type_cast_1355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1355_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1370_inst_req_0;
      type_cast_1370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1370_inst_req_1;
      type_cast_1370_inst_ack_1<= rack(0);
      type_cast_1370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp433_1367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv437_1371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack(0);
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr440_1377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv443_1381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1390_inst_req_0;
      type_cast_1390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1390_inst_req_1;
      type_cast_1390_inst_ack_1<= rack(0);
      type_cast_1390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr446_1387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv449_1391,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1400_inst_req_0;
      type_cast_1400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1400_inst_req_1;
      type_cast_1400_inst_ack_1<= rack(0);
      type_cast_1400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1400_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr452_1397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv455_1401,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1410_inst_req_0;
      type_cast_1410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1410_inst_req_1;
      type_cast_1410_inst_ack_1<= rack(0);
      type_cast_1410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr458_1407,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1420_inst_req_0;
      type_cast_1420_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1420_inst_req_1;
      type_cast_1420_inst_ack_1<= rack(0);
      type_cast_1420_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1420_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr464_1417,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv467_1421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1430_inst_req_0;
      type_cast_1430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1430_inst_req_1;
      type_cast_1430_inst_ack_1<= rack(0);
      type_cast_1430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr470_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv473_1431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1440_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1440_inst_req_0;
      type_cast_1440_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1440_inst_req_1;
      type_cast_1440_inst_ack_1<= rack(0);
      type_cast_1440_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1440_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr476_1437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1441,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_57,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_82,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_259_inst_req_0;
      type_cast_259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_259_inst_req_1;
      type_cast_259_inst_ack_1<= rack(0);
      type_cast_259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_289_inst_req_0;
      type_cast_289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_289_inst_req_1;
      type_cast_289_inst_ack_1<= rack(0);
      type_cast_289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_314_inst_req_0;
      type_cast_314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_314_inst_req_1;
      type_cast_314_inst_ack_1<= rack(0);
      type_cast_314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_327_inst_req_0;
      type_cast_327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_327_inst_req_1;
      type_cast_327_inst_ack_1<= rack(0);
      type_cast_327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_339_inst_req_0;
      type_cast_339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_339_inst_req_1;
      type_cast_339_inst_ack_1<= rack(0);
      type_cast_339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_352_inst_req_0;
      type_cast_352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_352_inst_req_1;
      type_cast_352_inst_ack_1<= rack(0);
      type_cast_352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_364_inst_req_0;
      type_cast_364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_364_inst_req_1;
      type_cast_364_inst_ack_1<= rack(0);
      type_cast_364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_377_inst_req_0;
      type_cast_377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_377_inst_req_1;
      type_cast_377_inst_ack_1<= rack(0);
      type_cast_377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_389_inst_req_0;
      type_cast_389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_389_inst_req_1;
      type_cast_389_inst_ack_1<= rack(0);
      type_cast_389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_402_inst_req_0;
      type_cast_402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_402_inst_req_1;
      type_cast_402_inst_ack_1<= rack(0);
      type_cast_402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp562x_xop_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_475_inst_req_0;
      type_cast_475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_475_inst_req_1;
      type_cast_475_inst_ack_1<= rack(0);
      type_cast_475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext556_626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_475_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_489_inst_req_0;
      type_cast_489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_489_inst_req_1;
      type_cast_489_inst_ack_1<= rack(0);
      type_cast_489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_502_inst_req_0;
      type_cast_502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_502_inst_req_1;
      type_cast_502_inst_ack_1<= rack(0);
      type_cast_502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_556_inst_req_0;
      type_cast_556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_556_inst_req_1;
      type_cast_556_inst_ack_1<= rack(0);
      type_cast_556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp548x_xop_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext540_833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_679_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_696_inst_req_0;
      type_cast_696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_696_inst_req_1;
      type_cast_696_inst_ack_1<= rack(0);
      type_cast_696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_693,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_745_inst_req_0;
      type_cast_745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_745_inst_req_1;
      type_cast_745_inst_ack_1<= rack(0);
      type_cast_745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_850_inst_req_0;
      type_cast_850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_850_inst_req_1;
      type_cast_850_inst_ack_1<= rack(0);
      type_cast_850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_858_inst_req_0;
      type_cast_858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_858_inst_req_1;
      type_cast_858_inst_ack_1<= rack(0);
      type_cast_858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp532x_xop_900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext526_945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_966_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1361_index_1_rename
    process(R_indvar_1360_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1360_resized;
      ov(13 downto 0) := iv;
      R_indvar_1360_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1361_index_1_resize
    process(indvar_1349) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1349;
      ov := iv(13 downto 0);
      R_indvar_1360_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1361_root_address_inst
    process(array_obj_ref_1361_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1361_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1361_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_rename
    process(R_indvar555_480_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar555_480_resized;
      ov(13 downto 0) := iv;
      R_indvar555_480_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_resize
    process(indvar555_469) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar555_469;
      ov := iv(13 downto 0);
      R_indvar555_480_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_root_address_inst
    process(array_obj_ref_481_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_481_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_481_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_rename
    process(R_indvar539_687_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar539_687_resized;
      ov(10 downto 0) := iv;
      R_indvar539_687_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_resize
    process(indvar539_676) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar539_676;
      ov := iv(10 downto 0);
      R_indvar539_687_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_root_address_inst
    process(array_obj_ref_688_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_688_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_rename
    process(R_indvar525_931_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar525_931_resized;
      ov(13 downto 0) := iv;
      R_indvar525_931_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_resize
    process(indvar525_920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar525_920;
      ov := iv(13 downto 0);
      R_indvar525_931_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_root_address_inst
    process(array_obj_ref_932_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_932_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_932_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1366_addr_0
    process(ptr_deref_1366_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1366_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1366_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1366_base_resize
    process(arrayidx432_1363) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx432_1363;
      ov := iv(13 downto 0);
      ptr_deref_1366_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1366_gather_scatter
    process(ptr_deref_1366_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1366_data_0;
      ov(63 downto 0) := iv;
      tmp433_1367 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1366_root_address_inst
    process(ptr_deref_1366_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1366_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1366_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_addr_0
    process(ptr_deref_618_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_base_resize
    process(arrayidx_483) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_483;
      ov := iv(13 downto 0);
      ptr_deref_618_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_gather_scatter
    process(add186_616) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_616;
      ov(63 downto 0) := iv;
      ptr_deref_618_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_root_address_inst
    process(ptr_deref_618_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_addr_0
    process(ptr_deref_825_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_base_resize
    process(arrayidx246_690) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_690;
      ov := iv(10 downto 0);
      ptr_deref_825_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_gather_scatter
    process(add242_823) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_823;
      ov(63 downto 0) := iv;
      ptr_deref_825_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_root_address_inst
    process(ptr_deref_825_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_addr_0
    process(ptr_deref_936_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_base_resize
    process(arrayidx269_934) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_934;
      ov := iv(13 downto 0);
      ptr_deref_936_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_gather_scatter
    process(type_cast_938_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_938_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_936_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_root_address_inst
    process(ptr_deref_936_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1305_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1305_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1305_branch_req_0,
          ack0 => if_stmt_1305_branch_ack_0,
          ack1 => if_stmt_1305_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1477_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1476;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1477_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1477_branch_req_0,
          ack0 => if_stmt_1477_branch_ack_0,
          ack1 => if_stmt_1477_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_416_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp513_415;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_416_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_416_branch_req_0,
          ack0 => if_stmt_416_branch_ack_0,
          ack1 => if_stmt_416_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_431_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194509_430;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_431_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_431_branch_req_0,
          ack0 => if_stmt_431_branch_ack_0,
          ack1 => if_stmt_431_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_632_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_631;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_632_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_632_branch_req_0,
          ack0 => if_stmt_632_branch_ack_0,
          ack1 => if_stmt_632_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_839_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_838;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_839_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_839_branch_req_0,
          ack0 => if_stmt_839_branch_ack_0,
          ack1 => if_stmt_839_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_876_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_876_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_876_branch_req_0,
          ack0 => if_stmt_876_branch_ack_0,
          ack1 => if_stmt_876_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_951_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_950;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_951_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_951_branch_req_0,
          ack0 => if_stmt_951_branch_ack_0,
          ack1 => if_stmt_951_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1328_inst
    process(tmp520_1317) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp520_1317, type_cast_1327_wire_constant, tmp_var);
      tmp520x_xop_1329 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_251_inst
    process(add74_247, shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_247, shr_235, tmp_var);
      add79_252 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_448_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_235, type_cast_447_wire_constant, tmp_var);
      tmp562x_xop_449 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_655_inst
    process(tmp548_644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp548_644, type_cast_654_wire_constant, tmp_var);
      tmp548x_xop_656 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_899_inst
    process(tmp532_888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp532_888, type_cast_898_wire_constant, tmp_var);
      tmp532x_xop_900 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1338_inst
    process(iNsTr_194_1333) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_194_1333, type_cast_1337_wire_constant, tmp_var);
      xx_xop_1339 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1470_inst
    process(indvar_1349) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1349, type_cast_1469_wire_constant, tmp_var);
      indvarx_xnext_1471 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_458_inst
    process(iNsTr_26_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_453, type_cast_457_wire_constant, tmp_var);
      xx_xop571_459 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_625_inst
    process(indvar555_469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar555_469, type_cast_624_wire_constant, tmp_var);
      indvarx_xnext556_626 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_665_inst
    process(iNsTr_39_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_660, type_cast_664_wire_constant, tmp_var);
      xx_xop570_666 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_832_inst
    process(indvar539_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar539_676, type_cast_831_wire_constant, tmp_var);
      indvarx_xnext540_833 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_909_inst
    process(iNsTr_53_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_904, type_cast_908_wire_constant, tmp_var);
      xx_xop569_910 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_944_inst
    process(indvar525_920) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar525_920, type_cast_943_wire_constant, tmp_var);
      indvarx_xnext526_945 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_246_inst
    process(iNsTr_14_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_241, type_cast_245_wire_constant, tmp_var);
      add74_247 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1475_inst
    process(indvarx_xnext_1471, tmp524_1346) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1471, tmp524_1346, tmp_var);
      exitcond1_1476 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_630_inst
    process(indvarx_xnext556_626, tmp567_466) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext556_626, tmp567_466, tmp_var);
      exitcond3_631 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_837_inst
    process(indvarx_xnext540_833, tmp553_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext540_833, tmp553_673, tmp_var);
      exitcond2_838 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_949_inst
    process(indvarx_xnext526_945, tmp537_917) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext526_945, tmp537_917, tmp_var);
      exitcond_950 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1044_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1043_wire_constant, tmp_var);
      shr304_1045 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1100_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1099_wire_constant, tmp_var);
      shr321_1101 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1156_inst
    process(add79_252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_252, type_cast_1155_wire_constant, tmp_var);
      shr338_1157 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1316_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_1315_wire_constant, tmp_var);
      tmp520_1317 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_234_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_233_wire_constant, tmp_var);
      shr_235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_239_wire_constant, tmp_var);
      iNsTr_14_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_643_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_283, type_cast_642_wire_constant, tmp_var);
      tmp548_644 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_887_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_886_wire_constant, tmp_var);
      tmp532_888 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1214_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1213_wire_constant, tmp_var);
      shr364_1215 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1224_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1223_wire_constant, tmp_var);
      shr370_1225 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1234_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1233_wire_constant, tmp_var);
      shr376_1235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1244_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1243_wire_constant, tmp_var);
      shr382_1245 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1254_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1253_wire_constant, tmp_var);
      shr388_1255 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1264_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1263_wire_constant, tmp_var);
      shr394_1265 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1274_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1273_wire_constant, tmp_var);
      shr400_1275 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1376_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1375_wire_constant, tmp_var);
      shr440_1377 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1386_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1385_wire_constant, tmp_var);
      shr446_1387 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1396_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1395_wire_constant, tmp_var);
      shr452_1397 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1406_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1405_wire_constant, tmp_var);
      shr458_1407 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1416_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1415_wire_constant, tmp_var);
      shr464_1417 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1426_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1425_wire_constant, tmp_var);
      shr470_1427 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1436_inst
    process(tmp433_1367) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1367, type_cast_1435_wire_constant, tmp_var);
      shr476_1437 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_223_inst
    process(conv63_215, conv61_211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_215, conv61_211, tmp_var);
      mul_224 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_228_inst
    process(mul_224, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_224, conv65_219, tmp_var);
      mul66_229 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_272_inst
    process(conv84_260, conv82_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_260, conv82_256, tmp_var);
      mul85_273 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_277_inst
    process(mul85_273, conv87_264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_273, conv87_264, tmp_var);
      mul88_278 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_282_inst
    process(mul88_278, conv90_268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_278, conv90_268, tmp_var);
      mul91_283 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_863_inst
    process(conv255_855, conv253_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_855, conv253_851, tmp_var);
      mul256_864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(mul256_864, conv258_859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_864, conv258_859, tmp_var);
      mul259_869 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_307_inst
    process(shl96_296, conv98_303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_296, conv98_303, tmp_var);
      add99_308 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_332_inst
    process(shl105_321, conv107_328) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_321, conv107_328, tmp_var);
      add108_333 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_357_inst
    process(shl114_346, conv116_353) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_346, conv116_353, tmp_var);
      add117_358 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_382_inst
    process(shl123_371, conv125_378) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_371, conv125_378, tmp_var);
      add126_383 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_407_inst
    process(shl132_396, conv134_403) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_396, conv134_403, tmp_var);
      add135_408 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_507_inst
    process(shl146_496, conv149_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_496, conv149_503, tmp_var);
      add150_508 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_525_inst
    process(shl152_514, conv155_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_514, conv155_521, tmp_var);
      add156_526 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_543_inst
    process(shl158_532, conv161_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_532, conv161_539, tmp_var);
      add162_544 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_561_inst
    process(shl164_550, conv167_557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_550, conv167_557, tmp_var);
      add168_562 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_579_inst
    process(shl170_568, conv173_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_568, conv173_575, tmp_var);
      add174_580 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_597_inst
    process(shl176_586, conv179_593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_586, conv179_593, tmp_var);
      add180_598 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_615_inst
    process(shl182_604, conv185_611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_604, conv185_611, tmp_var);
      add186_616 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_714_inst
    process(shl202_703, conv205_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_703, conv205_710, tmp_var);
      add206_715 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_732_inst
    process(shl208_721, conv211_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_721, conv211_728, tmp_var);
      add212_733 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_750_inst
    process(shl214_739, conv217_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_739, conv217_746, tmp_var);
      add218_751 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_768_inst
    process(shl220_757, conv223_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_757, conv223_764, tmp_var);
      add224_769 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_786_inst
    process(shl226_775, conv229_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_775, conv229_782, tmp_var);
      add230_787 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_804_inst
    process(shl232_793, conv235_800) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_793, conv235_800, tmp_var);
      add236_805 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_822_inst
    process(shl238_811, conv241_818) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_811, conv241_818, tmp_var);
      add242_823 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_295_inst
    process(conv95_290) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_290, type_cast_294_wire_constant, tmp_var);
      shl96_296 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_320_inst
    process(conv104_315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_315, type_cast_319_wire_constant, tmp_var);
      shl105_321 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_345_inst
    process(conv113_340) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_340, type_cast_344_wire_constant, tmp_var);
      shl114_346 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_370_inst
    process(conv122_365) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_365, type_cast_369_wire_constant, tmp_var);
      shl123_371 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_395_inst
    process(conv131_390) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_390, type_cast_394_wire_constant, tmp_var);
      shl132_396 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_495_inst
    process(conv144_490) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_490, type_cast_494_wire_constant, tmp_var);
      shl146_496 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_513_inst
    process(add150_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_508, type_cast_512_wire_constant, tmp_var);
      shl152_514 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_531_inst
    process(add156_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_526, type_cast_530_wire_constant, tmp_var);
      shl158_532 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_549_inst
    process(add162_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_544, type_cast_548_wire_constant, tmp_var);
      shl164_550 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_567_inst
    process(add168_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_562, type_cast_566_wire_constant, tmp_var);
      shl170_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_585_inst
    process(add174_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_580, type_cast_584_wire_constant, tmp_var);
      shl176_586 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_603_inst
    process(add180_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_598, type_cast_602_wire_constant, tmp_var);
      shl182_604 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_702_inst
    process(conv200_697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_697, type_cast_701_wire_constant, tmp_var);
      shl202_703 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_720_inst
    process(add206_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_715, type_cast_719_wire_constant, tmp_var);
      shl208_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_738_inst
    process(add212_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_733, type_cast_737_wire_constant, tmp_var);
      shl214_739 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_756_inst
    process(add218_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_751, type_cast_755_wire_constant, tmp_var);
      shl220_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_774_inst
    process(add224_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_769, type_cast_773_wire_constant, tmp_var);
      shl226_775 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_792_inst
    process(add230_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_787, type_cast_791_wire_constant, tmp_var);
      shl232_793 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_810_inst
    process(add236_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_805, type_cast_809_wire_constant, tmp_var);
      shl238_811 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1204_inst
    process(conv355_1200, conv276_968) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1200, conv276_968, tmp_var);
      sub_1205 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1322_inst
    process(tmp520_1317) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp520_1317, type_cast_1321_wire_constant, tmp_var);
      tmp521_1323 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_413_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_229, type_cast_412_wire_constant, tmp_var);
      cmp513_415 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_429_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_283, type_cast_428_wire_constant, tmp_var);
      cmp194509_430 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_442_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_235, type_cast_441_wire_constant, tmp_var);
      tmp563_443 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_649_inst
    process(tmp548_644) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp548_644, type_cast_648_wire_constant, tmp_var);
      tmp549_650 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_874_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_869, type_cast_873_wire_constant, tmp_var);
      cmp264505_875 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_893_inst
    process(tmp532_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp532_888, type_cast_892_wire_constant, tmp_var);
      tmp533_894 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1361_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1360_scaled;
      array_obj_ref_1361_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1361_index_offset_req_0;
      array_obj_ref_1361_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1361_index_offset_req_1;
      array_obj_ref_1361_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_481_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar555_480_scaled;
      array_obj_ref_481_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_481_index_offset_req_0;
      array_obj_ref_481_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_481_index_offset_req_1;
      array_obj_ref_481_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_688_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar539_687_scaled;
      array_obj_ref_688_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_688_index_offset_req_0;
      array_obj_ref_688_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_688_index_offset_req_1;
      array_obj_ref_688_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_932_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar525_931_scaled;
      array_obj_ref_932_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_932_index_offset_req_0;
      array_obj_ref_932_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_932_index_offset_req_1;
      array_obj_ref_932_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1198_inst
    process(call354_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1195, tmp_var);
      type_cast_1198_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_966_inst
    process(call275_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_962, tmp_var);
      type_cast_966_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1366_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1366_load_0_req_0;
      ptr_deref_1366_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1366_load_0_req_1;
      ptr_deref_1366_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1366_word_address_0;
      ptr_deref_1366_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_618_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_618_store_0_req_0;
      ptr_deref_618_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_618_store_0_req_1;
      ptr_deref_618_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_618_word_address_0;
      data_in <= ptr_deref_618_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_825_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_825_store_0_req_0;
      ptr_deref_825_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_825_store_0_req_1;
      ptr_deref_825_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_825_word_address_0;
      data_in <= ptr_deref_825_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_936_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_936_store_0_req_0;
      ptr_deref_936_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_936_store_0_req_1;
      ptr_deref_936_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_936_word_address_0;
      data_in <= ptr_deref_936_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1182_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1182_inst_req_0;
      RPIPE_Block0_done_1182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1182_inst_req_1;
      RPIPE_Block0_done_1182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1183 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1185_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1185_inst_req_0;
      RPIPE_Block1_done_1185_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1185_inst_req_1;
      RPIPE_Block1_done_1185_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1186 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1188_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1188_inst_req_0;
      RPIPE_Block2_done_1188_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1188_inst_req_1;
      RPIPE_Block2_done_1188_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1189 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1191_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1191_inst_req_0;
      RPIPE_Block3_done_1191_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1191_inst_req_1;
      RPIPE_Block3_done_1191_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1192 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_759_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_777_inst RPIPE_ConvTranspose_input_pipe_723_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_795_inst RPIPE_ConvTranspose_input_pipe_692_inst RPIPE_ConvTranspose_input_pipe_705_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_741_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_813_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_285_inst RPIPE_ConvTranspose_input_pipe_298_inst RPIPE_ConvTranspose_input_pipe_310_inst RPIPE_ConvTranspose_input_pipe_323_inst RPIPE_ConvTranspose_input_pipe_335_inst RPIPE_ConvTranspose_input_pipe_348_inst RPIPE_ConvTranspose_input_pipe_360_inst RPIPE_ConvTranspose_input_pipe_373_inst RPIPE_ConvTranspose_input_pipe_385_inst RPIPE_ConvTranspose_input_pipe_398_inst RPIPE_ConvTranspose_input_pipe_485_inst RPIPE_ConvTranspose_input_pipe_498_inst RPIPE_ConvTranspose_input_pipe_516_inst RPIPE_ConvTranspose_input_pipe_534_inst RPIPE_ConvTranspose_input_pipe_552_inst RPIPE_ConvTranspose_input_pipe_570_inst RPIPE_ConvTranspose_input_pipe_588_inst RPIPE_ConvTranspose_input_pipe_606_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call221_760 <= data_out(319 downto 312);
      call32_135 <= data_out(311 downto 304);
      call19_98 <= data_out(303 downto 296);
      call50_185 <= data_out(295 downto 288);
      call41_160 <= data_out(287 downto 280);
      call37_148 <= data_out(279 downto 272);
      call_35 <= data_out(271 downto 264);
      call5_60 <= data_out(263 downto 256);
      call46_173 <= data_out(255 downto 248);
      call227_778 <= data_out(247 downto 240);
      call209_724 <= data_out(239 downto 232);
      call23_110 <= data_out(231 downto 224);
      call28_123 <= data_out(223 downto 216);
      call14_85 <= data_out(215 downto 208);
      call233_796 <= data_out(207 downto 200);
      call199_693 <= data_out(199 downto 192);
      call203_706 <= data_out(191 downto 184);
      call2_48 <= data_out(183 downto 176);
      call215_742 <= data_out(175 downto 168);
      call10_73 <= data_out(167 downto 160);
      call239_814 <= data_out(159 downto 152);
      call55_198 <= data_out(151 downto 144);
      call92_286 <= data_out(143 downto 136);
      call97_299 <= data_out(135 downto 128);
      call101_311 <= data_out(127 downto 120);
      call106_324 <= data_out(119 downto 112);
      call110_336 <= data_out(111 downto 104);
      call115_349 <= data_out(103 downto 96);
      call119_361 <= data_out(95 downto 88);
      call124_374 <= data_out(87 downto 80);
      call128_386 <= data_out(79 downto 72);
      call133_399 <= data_out(71 downto 64);
      call143_486 <= data_out(63 downto 56);
      call147_499 <= data_out(55 downto 48);
      call153_517 <= data_out(47 downto 40);
      call159_535 <= data_out(39 downto 32);
      call165_553 <= data_out(31 downto 24);
      call171_571 <= data_out(23 downto 16);
      call177_589 <= data_out(15 downto 8);
      call183_607 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_993_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_996_inst WPIPE_Block0_start_1000_inst WPIPE_Block0_start_1004_inst WPIPE_Block0_start_1007_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_1010_inst WPIPE_Block0_start_969_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_972_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_981_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_996_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_1000_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_1004_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_1007_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_1010_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_969_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_972_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_981_inst_req_0;
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_996_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_1000_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_1004_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_1007_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_1010_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_969_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_972_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_996_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_1000_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_1004_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_1007_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_1010_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_969_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_972_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_981_inst_req_1;
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_996_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_1000_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_1004_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_1007_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_1010_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_969_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_972_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_333 & add99_308 & type_cast_998_wire_constant & type_cast_1002_wire_constant & add117_358 & add126_383 & add48_182 & add135_408 & add_57 & add57_207 & add12_82 & add21_107 & add30_132 & add39_157;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1063_inst WPIPE_Block1_start_1060_inst WPIPE_Block1_start_1050_inst WPIPE_Block1_start_1066_inst WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1034_inst WPIPE_Block1_start_1037_inst WPIPE_Block1_start_1057_inst WPIPE_Block1_start_1013_inst WPIPE_Block1_start_1016_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1028_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1063_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1060_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1050_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1037_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1057_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1013_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1016_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1028_inst_req_0;
      WPIPE_Block1_start_1063_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1060_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1050_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1057_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1013_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1016_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1063_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1060_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1050_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1034_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1037_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1057_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1013_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1016_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1028_inst_req_1;
      WPIPE_Block1_start_1063_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1060_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1050_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1034_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1057_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1013_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1016_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_383 & add117_358 & conv305_1049 & add135_408 & add57_207 & add99_308 & add108_333 & conv307_1056 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1116_inst WPIPE_Block2_start_1122_inst WPIPE_Block2_start_1069_inst WPIPE_Block2_start_1072_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1090_inst WPIPE_Block2_start_1093_inst WPIPE_Block2_start_1106_inst WPIPE_Block2_start_1113_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1116_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1122_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1069_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1072_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1090_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1093_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1106_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1113_inst_req_0;
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1116_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1069_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1072_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1090_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1093_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1106_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1113_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1116_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1122_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1069_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1072_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1090_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1093_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1106_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1113_inst_req_1;
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1116_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1069_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1072_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1090_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1093_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1106_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1113_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_383 & add117_358 & add135_408 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308 & add108_333 & conv322_1105 & conv324_1112;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1149_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1162_inst WPIPE_Block3_start_1172_inst WPIPE_Block3_start_1175_inst WPIPE_Block3_start_1146_inst WPIPE_Block3_start_1128_inst WPIPE_Block3_start_1143_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1125_inst WPIPE_Block3_start_1169_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1162_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1172_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1175_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1146_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1128_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1143_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1125_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1169_inst_req_0;
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1162_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1172_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1146_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1128_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1125_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1169_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1149_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1162_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1172_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1175_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1146_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1128_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1143_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1125_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1169_inst_req_1;
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1149_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1162_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1172_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1146_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1128_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1125_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1169_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add39_157 & add108_333 & add48_182 & add21_107 & add30_132 & conv339_1161 & add117_358 & add126_383 & add99_308 & add12_82 & add57_207 & add135_408 & add_57 & conv341_1168;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1292_inst WPIPE_ConvTranspose_output_pipe_1295_inst WPIPE_ConvTranspose_output_pipe_1280_inst WPIPE_ConvTranspose_output_pipe_1289_inst WPIPE_ConvTranspose_output_pipe_1283_inst WPIPE_ConvTranspose_output_pipe_1286_inst WPIPE_ConvTranspose_output_pipe_1301_inst WPIPE_ConvTranspose_output_pipe_1298_inst WPIPE_ConvTranspose_output_pipe_1442_inst WPIPE_ConvTranspose_output_pipe_1445_inst WPIPE_ConvTranspose_output_pipe_1448_inst WPIPE_ConvTranspose_output_pipe_1451_inst WPIPE_ConvTranspose_output_pipe_1454_inst WPIPE_ConvTranspose_output_pipe_1457_inst WPIPE_ConvTranspose_output_pipe_1460_inst WPIPE_ConvTranspose_output_pipe_1463_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1457_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1460_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1463_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1457_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1460_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1463_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv379_1239 & conv373_1229 & conv403_1279 & conv385_1249 & conv397_1269 & conv391_1259 & conv361_1209 & conv367_1219 & conv479_1441 & conv473_1431 & conv467_1421 & conv461_1411 & conv455_1401 & conv449_1391 & conv443_1381 & conv437_1371;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1195_call call_stmt_962_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1195_call_req_0;
      reqL_unguarded(0) <= call_stmt_962_call_req_0;
      call_stmt_1195_call_ack_0 <= ackL_unguarded(1);
      call_stmt_962_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1195_call_req_1;
      reqR_unguarded(0) <= call_stmt_962_call_req_1;
      call_stmt_1195_call_ack_1 <= ackR_unguarded(1);
      call_stmt_962_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call354_1195 <= data_out(127 downto 64);
      call275_962 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3758_start: Boolean;
  signal convTransposeA_CP_3758_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1600_ack_0 : boolean;
  signal type_cast_1821_inst_ack_1 : boolean;
  signal type_cast_1827_inst_ack_1 : boolean;
  signal type_cast_1827_inst_req_1 : boolean;
  signal phi_stmt_1822_req_1 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal phi_stmt_1614_req_0 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal type_cast_1819_inst_ack_0 : boolean;
  signal type_cast_1819_inst_req_1 : boolean;
  signal phi_stmt_1614_ack_0 : boolean;
  signal phi_stmt_1816_req_1 : boolean;
  signal type_cast_1815_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1819_inst_ack_1 : boolean;
  signal phi_stmt_1607_ack_0 : boolean;
  signal phi_stmt_1816_req_0 : boolean;
  signal type_cast_1815_inst_ack_0 : boolean;
  signal phi_stmt_1822_ack_0 : boolean;
  signal phi_stmt_1621_ack_0 : boolean;
  signal type_cast_1821_inst_req_1 : boolean;
  signal type_cast_1819_inst_req_0 : boolean;
  signal phi_stmt_1621_req_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1496_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1514_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1514_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1505_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1505_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1496_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1508_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1508_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1496_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1502_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1502_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1496_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1508_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1508_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1502_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1505_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1505_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1502_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1511_inst_req_1 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1514_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1514_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1517_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1517_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1517_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1517_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1520_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1520_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1520_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1520_inst_ack_1 : boolean;
  signal type_cast_1524_inst_req_0 : boolean;
  signal type_cast_1524_inst_ack_0 : boolean;
  signal type_cast_1524_inst_req_1 : boolean;
  signal type_cast_1524_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1533_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1533_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1533_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1533_inst_ack_1 : boolean;
  signal type_cast_1537_inst_req_0 : boolean;
  signal type_cast_1537_inst_ack_0 : boolean;
  signal type_cast_1537_inst_req_1 : boolean;
  signal type_cast_1537_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1545_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1545_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1545_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1545_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1548_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1548_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1548_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1548_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1551_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1551_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1551_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1551_inst_ack_1 : boolean;
  signal type_cast_1578_inst_req_0 : boolean;
  signal type_cast_1578_inst_ack_0 : boolean;
  signal type_cast_1578_inst_req_1 : boolean;
  signal type_cast_1578_inst_ack_1 : boolean;
  signal type_cast_1582_inst_req_0 : boolean;
  signal type_cast_1582_inst_ack_0 : boolean;
  signal type_cast_1582_inst_req_1 : boolean;
  signal type_cast_1582_inst_ack_1 : boolean;
  signal type_cast_1586_inst_req_0 : boolean;
  signal type_cast_1586_inst_ack_0 : boolean;
  signal type_cast_1586_inst_req_1 : boolean;
  signal type_cast_1586_inst_ack_1 : boolean;
  signal type_cast_1590_inst_req_0 : boolean;
  signal type_cast_1590_inst_ack_0 : boolean;
  signal type_cast_1590_inst_req_1 : boolean;
  signal type_cast_1590_inst_ack_1 : boolean;
  signal type_cast_1662_inst_req_0 : boolean;
  signal type_cast_1662_inst_ack_0 : boolean;
  signal type_cast_1662_inst_req_1 : boolean;
  signal type_cast_1662_inst_ack_1 : boolean;
  signal type_cast_1666_inst_req_0 : boolean;
  signal type_cast_1666_inst_ack_0 : boolean;
  signal type_cast_1666_inst_req_1 : boolean;
  signal type_cast_1666_inst_ack_1 : boolean;
  signal type_cast_1670_inst_req_0 : boolean;
  signal type_cast_1670_inst_ack_0 : boolean;
  signal type_cast_1670_inst_req_1 : boolean;
  signal type_cast_1670_inst_ack_1 : boolean;
  signal type_cast_1700_inst_req_0 : boolean;
  signal type_cast_1700_inst_ack_0 : boolean;
  signal type_cast_1700_inst_req_1 : boolean;
  signal type_cast_1700_inst_ack_1 : boolean;
  signal phi_stmt_1621_req_1 : boolean;
  signal type_cast_1627_inst_ack_1 : boolean;
  signal type_cast_1627_inst_req_1 : boolean;
  signal phi_stmt_1816_ack_0 : boolean;
  signal array_obj_ref_1706_index_offset_req_0 : boolean;
  signal array_obj_ref_1706_index_offset_ack_0 : boolean;
  signal array_obj_ref_1706_index_offset_req_1 : boolean;
  signal array_obj_ref_1706_index_offset_ack_1 : boolean;
  signal phi_stmt_1809_ack_0 : boolean;
  signal addr_of_1707_final_reg_req_0 : boolean;
  signal addr_of_1707_final_reg_ack_0 : boolean;
  signal addr_of_1707_final_reg_req_1 : boolean;
  signal addr_of_1707_final_reg_ack_1 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal type_cast_1827_inst_ack_0 : boolean;
  signal type_cast_1827_inst_req_0 : boolean;
  signal type_cast_1627_inst_ack_0 : boolean;
  signal type_cast_1627_inst_req_0 : boolean;
  signal ptr_deref_1711_load_0_req_0 : boolean;
  signal ptr_deref_1711_load_0_ack_0 : boolean;
  signal phi_stmt_1607_req_1 : boolean;
  signal ptr_deref_1711_load_0_req_1 : boolean;
  signal ptr_deref_1711_load_0_ack_1 : boolean;
  signal phi_stmt_1809_req_0 : boolean;
  signal phi_stmt_1822_req_0 : boolean;
  signal array_obj_ref_1729_index_offset_req_0 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal array_obj_ref_1729_index_offset_ack_0 : boolean;
  signal array_obj_ref_1729_index_offset_req_1 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal array_obj_ref_1729_index_offset_ack_1 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal phi_stmt_1809_req_1 : boolean;
  signal type_cast_1815_inst_ack_1 : boolean;
  signal type_cast_1815_inst_req_1 : boolean;
  signal addr_of_1730_final_reg_req_0 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal addr_of_1730_final_reg_ack_0 : boolean;
  signal addr_of_1730_final_reg_req_1 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal addr_of_1730_final_reg_ack_1 : boolean;
  signal phi_stmt_1614_req_1 : boolean;
  signal type_cast_1620_inst_ack_1 : boolean;
  signal type_cast_1620_inst_req_1 : boolean;
  signal type_cast_1620_inst_ack_0 : boolean;
  signal type_cast_1620_inst_req_0 : boolean;
  signal phi_stmt_1600_req_1 : boolean;
  signal ptr_deref_1733_store_0_req_0 : boolean;
  signal ptr_deref_1733_store_0_ack_0 : boolean;
  signal ptr_deref_1733_store_0_req_1 : boolean;
  signal ptr_deref_1733_store_0_ack_1 : boolean;
  signal type_cast_1738_inst_req_0 : boolean;
  signal type_cast_1738_inst_ack_0 : boolean;
  signal type_cast_1738_inst_req_1 : boolean;
  signal type_cast_1738_inst_ack_1 : boolean;
  signal if_stmt_1751_branch_req_0 : boolean;
  signal if_stmt_1751_branch_ack_1 : boolean;
  signal if_stmt_1751_branch_ack_0 : boolean;
  signal type_cast_1779_inst_req_0 : boolean;
  signal type_cast_1779_inst_ack_0 : boolean;
  signal type_cast_1779_inst_req_1 : boolean;
  signal type_cast_1779_inst_ack_1 : boolean;
  signal type_cast_1795_inst_req_0 : boolean;
  signal type_cast_1795_inst_ack_0 : boolean;
  signal type_cast_1795_inst_req_1 : boolean;
  signal type_cast_1795_inst_ack_1 : boolean;
  signal if_stmt_1802_branch_req_0 : boolean;
  signal if_stmt_1802_branch_ack_1 : boolean;
  signal if_stmt_1802_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1838_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1838_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1838_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1838_inst_ack_1 : boolean;
  signal phi_stmt_1600_req_0 : boolean;
  signal phi_stmt_1607_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3758_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3758: Block -- control-path 
    signal convTransposeA_CP_3758_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3758_elements(0) <= convTransposeA_CP_3758_start;
    convTransposeA_CP_3758_symbol <= convTransposeA_CP_3758_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1491/branch_block_stmt_1491__entry__
      -- CP-element group 0: 	 branch_block_stmt_1491/$entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552__entry__
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/$entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Update/cr
      -- 
    rr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => RPIPE_Block0_start_1493_inst_req_0); -- 
    cr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => type_cast_1524_inst_req_1); -- 
    cr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => type_cast_1537_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/merge_stmt_1808__exit__
      -- CP-element group 1: 	 branch_block_stmt_1491/assign_stmt_1834__entry__
      -- CP-element group 1: 	 branch_block_stmt_1491/assign_stmt_1834__exit__
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/assign_stmt_1834/$entry
      -- CP-element group 1: 	 branch_block_stmt_1491/assign_stmt_1834/$exit
      -- 
    rr_4515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1613_inst_req_0); -- 
    cr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1613_inst_req_1); -- 
    cr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1606_inst_req_1); -- 
    cr_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1627_inst_req_1); -- 
    rr_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1606_inst_req_0); -- 
    rr_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1627_inst_req_0); -- 
    cr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1620_inst_req_1); -- 
    rr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1620_inst_req_0); -- 
    convTransposeA_CP_3758_elements(1) <= convTransposeA_CP_3758_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Update/cr
      -- 
    ra_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1493_inst_ack_0, ack => convTransposeA_CP_3758_elements(2)); -- 
    cr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(2), ack => RPIPE_Block0_start_1493_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1493_Update/$exit
      -- 
    ca_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1493_inst_ack_1, ack => convTransposeA_CP_3758_elements(3)); -- 
    rr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(3), ack => RPIPE_Block0_start_1496_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Update/cr
      -- 
    ra_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1496_inst_ack_0, ack => convTransposeA_CP_3758_elements(4)); -- 
    cr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(4), ack => RPIPE_Block0_start_1496_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1496_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_sample_start_
      -- 
    ca_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1496_inst_ack_1, ack => convTransposeA_CP_3758_elements(5)); -- 
    rr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(5), ack => RPIPE_Block0_start_1499_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_sample_completed_
      -- 
    ra_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_0, ack => convTransposeA_CP_3758_elements(6)); -- 
    cr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(6), ack => RPIPE_Block0_start_1499_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1499_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Sample/rr
      -- 
    ca_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_1, ack => convTransposeA_CP_3758_elements(7)); -- 
    rr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(7), ack => RPIPE_Block0_start_1502_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Update/cr
      -- 
    ra_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1502_inst_ack_0, ack => convTransposeA_CP_3758_elements(8)); -- 
    cr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(8), ack => RPIPE_Block0_start_1502_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1502_Update/ca
      -- 
    ca_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1502_inst_ack_1, ack => convTransposeA_CP_3758_elements(9)); -- 
    rr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(9), ack => RPIPE_Block0_start_1505_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Sample/ra
      -- 
    ra_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1505_inst_ack_0, ack => convTransposeA_CP_3758_elements(10)); -- 
    cr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(10), ack => RPIPE_Block0_start_1505_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1505_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Sample/rr
      -- 
    ca_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1505_inst_ack_1, ack => convTransposeA_CP_3758_elements(11)); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(11), ack => RPIPE_Block0_start_1508_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Sample/ra
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1508_inst_ack_0, ack => convTransposeA_CP_3758_elements(12)); -- 
    cr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(12), ack => RPIPE_Block0_start_1508_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1508_Update/$exit
      -- 
    ca_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1508_inst_ack_1, ack => convTransposeA_CP_3758_elements(13)); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(13), ack => RPIPE_Block0_start_1511_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Update/cr
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1511_inst_ack_0, ack => convTransposeA_CP_3758_elements(14)); -- 
    cr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(14), ack => RPIPE_Block0_start_1511_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1511_Update/$exit
      -- 
    ca_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1511_inst_ack_1, ack => convTransposeA_CP_3758_elements(15)); -- 
    rr_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(15), ack => RPIPE_Block0_start_1514_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Update/cr
      -- 
    ra_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1514_inst_ack_0, ack => convTransposeA_CP_3758_elements(16)); -- 
    cr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(16), ack => RPIPE_Block0_start_1514_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1514_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Sample/rr
      -- 
    ca_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1514_inst_ack_1, ack => convTransposeA_CP_3758_elements(17)); -- 
    rr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(17), ack => RPIPE_Block0_start_1517_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Update/cr
      -- 
    ra_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1517_inst_ack_0, ack => convTransposeA_CP_3758_elements(18)); -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(18), ack => RPIPE_Block0_start_1517_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1517_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Sample/rr
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1517_inst_ack_1, ack => convTransposeA_CP_3758_elements(19)); -- 
    rr_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(19), ack => RPIPE_Block0_start_1520_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Update/cr
      -- 
    ra_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1520_inst_ack_0, ack => convTransposeA_CP_3758_elements(20)); -- 
    cr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(20), ack => RPIPE_Block0_start_1520_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1520_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Sample/rr
      -- 
    ca_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1520_inst_ack_1, ack => convTransposeA_CP_3758_elements(21)); -- 
    rr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(21), ack => type_cast_1524_inst_req_0); -- 
    rr_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(21), ack => RPIPE_Block0_start_1533_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Sample/ra
      -- 
    ra_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1524_inst_ack_0, ack => convTransposeA_CP_3758_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1524_Update/ca
      -- 
    ca_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1524_inst_ack_1, ack => convTransposeA_CP_3758_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Update/cr
      -- 
    ra_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1533_inst_ack_0, ack => convTransposeA_CP_3758_elements(24)); -- 
    cr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(24), ack => RPIPE_Block0_start_1533_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1533_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Sample/rr
      -- 
    ca_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1533_inst_ack_1, ack => convTransposeA_CP_3758_elements(25)); -- 
    rr_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(25), ack => type_cast_1537_inst_req_0); -- 
    rr_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(25), ack => RPIPE_Block0_start_1545_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Sample/ra
      -- 
    ra_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1537_inst_ack_0, ack => convTransposeA_CP_3758_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/type_cast_1537_Update/ca
      -- 
    ca_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1537_inst_ack_1, ack => convTransposeA_CP_3758_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Update/cr
      -- 
    ra_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1545_inst_ack_0, ack => convTransposeA_CP_3758_elements(28)); -- 
    cr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(28), ack => RPIPE_Block0_start_1545_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1545_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Sample/rr
      -- 
    ca_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1545_inst_ack_1, ack => convTransposeA_CP_3758_elements(29)); -- 
    rr_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(29), ack => RPIPE_Block0_start_1548_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Update/cr
      -- 
    ra_4003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1548_inst_ack_0, ack => convTransposeA_CP_3758_elements(30)); -- 
    cr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(30), ack => RPIPE_Block0_start_1548_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1548_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Sample/rr
      -- 
    ca_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1548_inst_ack_1, ack => convTransposeA_CP_3758_elements(31)); -- 
    rr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(31), ack => RPIPE_Block0_start_1551_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Update/cr
      -- 
    ra_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1551_inst_ack_0, ack => convTransposeA_CP_3758_elements(32)); -- 
    cr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(32), ack => RPIPE_Block0_start_1551_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/RPIPE_Block0_start_1551_Update/ca
      -- 
    ca_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1551_inst_ack_1, ack => convTransposeA_CP_3758_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552__exit__
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1494_to_assign_stmt_1552/$exit
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597__entry__
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Update/cr
      -- 
    rr_4033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1578_inst_req_0); -- 
    cr_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1578_inst_req_1); -- 
    rr_4047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1582_inst_req_0); -- 
    cr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1582_inst_req_1); -- 
    rr_4061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1586_inst_req_0); -- 
    cr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1586_inst_req_1); -- 
    rr_4075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1590_inst_req_0); -- 
    cr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1590_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(23) & convTransposeA_CP_3758_elements(27) & convTransposeA_CP_3758_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Sample/ra
      -- 
    ra_4034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1578_inst_ack_0, ack => convTransposeA_CP_3758_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1578_Update/ca
      -- 
    ca_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1578_inst_ack_1, ack => convTransposeA_CP_3758_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Sample/ra
      -- 
    ra_4048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1582_inst_ack_0, ack => convTransposeA_CP_3758_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1582_Update/ca
      -- 
    ca_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1582_inst_ack_1, ack => convTransposeA_CP_3758_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Sample/ra
      -- 
    ra_4062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1586_inst_ack_0, ack => convTransposeA_CP_3758_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1586_Update/ca
      -- 
    ca_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1586_inst_ack_1, ack => convTransposeA_CP_3758_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Sample/ra
      -- 
    ra_4076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_0, ack => convTransposeA_CP_3758_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/type_cast_1590_Update/ca
      -- 
    ca_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_1, ack => convTransposeA_CP_3758_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597__exit__
      -- CP-element group 43: 	 branch_block_stmt_1491/assign_stmt_1559_to_assign_stmt_1597/$exit
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/$entry
      -- CP-element group 43: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(36) & convTransposeA_CP_3758_elements(38) & convTransposeA_CP_3758_elements(40) & convTransposeA_CP_3758_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Sample/ra
      -- 
    ra_4093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_0, ack => convTransposeA_CP_3758_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Update/ca
      -- 
    ca_4098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_1, ack => convTransposeA_CP_3758_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Sample/ra
      -- 
    ra_4107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_0, ack => convTransposeA_CP_3758_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Update/ca
      -- 
    ca_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1666_inst_ack_1, ack => convTransposeA_CP_3758_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Sample/ra
      -- 
    ra_4121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_0, ack => convTransposeA_CP_3758_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Update/ca
      -- 
    ca_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_1, ack => convTransposeA_CP_3758_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Sample/ra
      -- 
    ra_4135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1700_inst_ack_0, ack => convTransposeA_CP_3758_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Sample/req
      -- 
    ca_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1700_inst_ack_1, ack => convTransposeA_CP_3758_elements(51)); -- 
    req_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(51), ack => array_obj_ref_1706_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Sample/ack
      -- 
    ack_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1706_index_offset_ack_0, ack => convTransposeA_CP_3758_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_request/req
      -- 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1706_index_offset_ack_1, ack => convTransposeA_CP_3758_elements(53)); -- 
    req_4180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(53), ack => addr_of_1707_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_request/ack
      -- 
    ack_4181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1707_final_reg_ack_0, ack => convTransposeA_CP_3758_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/word_0/rr
      -- 
    ack_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1707_final_reg_ack_1, ack => convTransposeA_CP_3758_elements(55)); -- 
    rr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(55), ack => ptr_deref_1711_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Sample/word_access_start/word_0/ra
      -- 
    ra_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1711_load_0_ack_0, ack => convTransposeA_CP_3758_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/ptr_deref_1711_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/ptr_deref_1711_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/ptr_deref_1711_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/ptr_deref_1711_Merge/merge_ack
      -- 
    ca_4231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1711_load_0_ack_1, ack => convTransposeA_CP_3758_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Sample/req
      -- 
    req_4261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(58), ack => array_obj_ref_1729_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(45) & convTransposeA_CP_3758_elements(47) & convTransposeA_CP_3758_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Sample/ack
      -- 
    ack_4262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1729_index_offset_ack_0, ack => convTransposeA_CP_3758_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_request/req
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1729_index_offset_ack_1, ack => convTransposeA_CP_3758_elements(60)); -- 
    req_4276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(60), ack => addr_of_1730_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_request/ack
      -- 
    ack_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1730_final_reg_ack_0, ack => convTransposeA_CP_3758_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_word_addrgen/root_register_ack
      -- 
    ack_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1730_final_reg_ack_1, ack => convTransposeA_CP_3758_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/ptr_deref_1733_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/ptr_deref_1733_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/ptr_deref_1733_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/ptr_deref_1733_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/word_0/rr
      -- 
    rr_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(63), ack => ptr_deref_1733_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(57) & convTransposeA_CP_3758_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Sample/word_access_start/word_0/ra
      -- 
    ra_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1733_store_0_ack_0, ack => convTransposeA_CP_3758_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/word_0/ca
      -- 
    ca_4332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1733_store_0_ack_1, ack => convTransposeA_CP_3758_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Sample/ra
      -- 
    ra_4341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_0, ack => convTransposeA_CP_3758_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Update/ca
      -- 
    ca_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_1, ack => convTransposeA_CP_3758_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751__entry__
      -- CP-element group 68: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750__exit__
      -- CP-element group 68: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/$exit
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1491/R_cmp_1752_place
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1491/if_stmt_1751_else_link/$entry
      -- 
    branch_req_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(68), ack => if_stmt_1751_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(52) & convTransposeA_CP_3758_elements(59) & convTransposeA_CP_3758_elements(65) & convTransposeA_CP_3758_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1491/merge_stmt_1757_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/merge_stmt_1757_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1491/merge_stmt_1757_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/merge_stmt_1757_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1491/merge_stmt_1757__exit__
      -- CP-element group 69: 	 branch_block_stmt_1491/assign_stmt_1763__entry__
      -- CP-element group 69: 	 branch_block_stmt_1491/assign_stmt_1763__exit__
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1491/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/if_stmt_1751_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1491/if_stmt_1751_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1491/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1491/assign_stmt_1763/$entry
      -- CP-element group 69: 	 branch_block_stmt_1491/assign_stmt_1763/$exit
      -- 
    if_choice_transition_4359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1751_branch_ack_1, ack => convTransposeA_CP_3758_elements(69)); -- 
    cr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1827_inst_req_1); -- 
    rr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1815_inst_req_0); -- 
    cr_4704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1821_inst_req_1); -- 
    rr_4699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1821_inst_req_0); -- 
    rr_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1827_inst_req_0); -- 
    cr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1815_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1491/merge_stmt_1765_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1491/merge_stmt_1765_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1491/merge_stmt_1765_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1491/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/merge_stmt_1765_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801__entry__
      -- CP-element group 70: 	 branch_block_stmt_1491/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1491/merge_stmt_1765__exit__
      -- CP-element group 70: 	 branch_block_stmt_1491/if_stmt_1751_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1491/if_stmt_1751_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1491/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Update/cr
      -- 
    else_choice_transition_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1751_branch_ack_0, ack => convTransposeA_CP_3758_elements(70)); -- 
    rr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1779_inst_req_0); -- 
    cr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1779_inst_req_1); -- 
    cr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1795_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Sample/ra
      -- 
    ra_4380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_0, ack => convTransposeA_CP_3758_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1779_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Sample/rr
      -- 
    ca_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1779_inst_ack_1, ack => convTransposeA_CP_3758_elements(72)); -- 
    rr_4393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(72), ack => type_cast_1795_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Sample/ra
      -- 
    ra_4394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_0, ack => convTransposeA_CP_3758_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801__exit__
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802__entry__
      -- CP-element group 74: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/$exit
      -- CP-element group 74: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1491/assign_stmt_1771_to_assign_stmt_1801/type_cast_1795_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1491/R_cmp112_1803_place
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1491/if_stmt_1802_else_link/$entry
      -- 
    ca_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_1, ack => convTransposeA_CP_3758_elements(74)); -- 
    branch_req_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(74), ack => if_stmt_1802_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1491/merge_stmt_1836_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1491/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1491/merge_stmt_1836__exit__
      -- CP-element group 75: 	 branch_block_stmt_1491/assign_stmt_1841__entry__
      -- CP-element group 75: 	 branch_block_stmt_1491/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1491/merge_stmt_1836_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1491/merge_stmt_1836_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1491/merge_stmt_1836_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1491/if_stmt_1802_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1491/if_stmt_1802_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1491/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1491/assign_stmt_1841/$entry
      -- CP-element group 75: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Sample/req
      -- 
    if_choice_transition_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1802_branch_ack_1, ack => convTransposeA_CP_3758_elements(75)); -- 
    req_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(75), ack => WPIPE_Block0_done_1838_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1491/if_stmt_1802_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1491/if_stmt_1802_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1802_branch_ack_0, ack => convTransposeA_CP_3758_elements(76)); -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1819_inst_req_1); -- 
    rr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1819_inst_req_0); -- 
    cr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1825_inst_req_1); -- 
    rr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1825_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Update/req
      -- 
    ack_4433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1838_inst_ack_0, ack => convTransposeA_CP_3758_elements(77)); -- 
    req_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(77), ack => WPIPE_Block0_done_1838_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1491/merge_stmt_1843_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1491/merge_stmt_1843_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1491/assign_stmt_1841__exit__
      -- CP-element group 78: 	 branch_block_stmt_1491/merge_stmt_1843_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1491/merge_stmt_1843_PhiAck/dummy
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1491/branch_block_stmt_1491__exit__
      -- CP-element group 78: 	 branch_block_stmt_1491/merge_stmt_1843__exit__
      -- CP-element group 78: 	 branch_block_stmt_1491/$exit
      -- CP-element group 78: 	 branch_block_stmt_1491/return__
      -- CP-element group 78: 	 branch_block_stmt_1491/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1491/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1491/assign_stmt_1841/$exit
      -- CP-element group 78: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1491/assign_stmt_1841/WPIPE_Block0_done_1838_Update/ack
      -- 
    ack_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1838_inst_ack_1, ack => convTransposeA_CP_3758_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/$exit
      -- CP-element group 79: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1604_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_req
      -- 
    phi_stmt_1600_req_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1600_req_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(79), ack => phi_stmt_1600_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/$exit
      -- CP-element group 80: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1611_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_req
      -- 
    phi_stmt_1607_req_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1607_req_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(80), ack => phi_stmt_1607_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_req
      -- CP-element group 81: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1618_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1614/$exit
      -- 
    phi_stmt_1614_req_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1614_req_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(81), ack => phi_stmt_1614_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/$exit
      -- CP-element group 82: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1625_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- 
    phi_stmt_1621_req_4473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(82), ack => phi_stmt_1621_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1491/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(79) & convTransposeA_CP_3758_elements(80) & convTransposeA_CP_3758_elements(81) & convTransposeA_CP_3758_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Sample/$exit
      -- 
    ra_4493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => convTransposeA_CP_3758_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/Update/$exit
      -- 
    ca_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => convTransposeA_CP_3758_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/$exit
      -- CP-element group 86: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/$exit
      -- CP-element group 86: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_sources/type_cast_1606/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1600/phi_stmt_1600_req
      -- 
    phi_stmt_1600_req_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1600_req_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(86), ack => phi_stmt_1600_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(84) & convTransposeA_CP_3758_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Sample/ra
      -- 
    ra_4516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => convTransposeA_CP_3758_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/Update/ca
      -- 
    ca_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => convTransposeA_CP_3758_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_req
      -- CP-element group 89: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/type_cast_1613/$exit
      -- CP-element group 89: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/phi_stmt_1607_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1607/$exit
      -- 
    phi_stmt_1607_req_4522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1607_req_4522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(89), ack => phi_stmt_1607_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(87) & convTransposeA_CP_3758_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Sample/ra
      -- 
    ra_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_0, ack => convTransposeA_CP_3758_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/Update/$exit
      -- 
    ca_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1620_inst_ack_1, ack => convTransposeA_CP_3758_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/$exit
      -- CP-element group 92: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/type_cast_1620/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/$exit
      -- CP-element group 92: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1614/phi_stmt_1614_req
      -- 
    phi_stmt_1614_req_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1614_req_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(92), ack => phi_stmt_1614_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(90) & convTransposeA_CP_3758_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Sample/$exit
      -- 
    ra_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_0, ack => convTransposeA_CP_3758_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/Update/$exit
      -- 
    ca_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1627_inst_ack_1, ack => convTransposeA_CP_3758_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_req
      -- CP-element group 95: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/type_cast_1627/$exit
      -- CP-element group 95: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/phi_stmt_1621_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1621/$exit
      -- 
    phi_stmt_1621_req_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1621_req_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(95), ack => phi_stmt_1621_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(93) & convTransposeA_CP_3758_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1491/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(86) & convTransposeA_CP_3758_elements(89) & convTransposeA_CP_3758_elements(92) & convTransposeA_CP_3758_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/$entry
      -- CP-element group 97: 	 branch_block_stmt_1491/merge_stmt_1599_PhiReqMerge
      -- 
    convTransposeA_CP_3758_elements(97) <= OrReduce(convTransposeA_CP_3758_elements(83) & convTransposeA_CP_3758_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/phi_stmt_1600_ack
      -- 
    phi_stmt_1600_ack_4573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1600_ack_0, ack => convTransposeA_CP_3758_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/phi_stmt_1607_ack
      -- 
    phi_stmt_1607_ack_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1607_ack_0, ack => convTransposeA_CP_3758_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/phi_stmt_1614_ack
      -- 
    phi_stmt_1614_ack_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1614_ack_0, ack => convTransposeA_CP_3758_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/phi_stmt_1621_ack
      -- 
    phi_stmt_1621_ack_4576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1621_ack_0, ack => convTransposeA_CP_3758_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1491/merge_stmt_1599_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1491/merge_stmt_1599__exit__
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750__entry__
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1662_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1666_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1670_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1700_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1706_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1707_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1711_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/array_obj_ref_1729_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/addr_of_1730_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/ptr_deref_1733_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1491/assign_stmt_1634_to_assign_stmt_1750/type_cast_1738_Update/cr
      -- 
    rr_4092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1662_inst_req_0); -- 
    cr_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1662_inst_req_1); -- 
    rr_4106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1666_inst_req_0); -- 
    cr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1666_inst_req_1); -- 
    rr_4120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1670_inst_req_0); -- 
    cr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1670_inst_req_1); -- 
    rr_4134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1700_inst_req_0); -- 
    cr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1700_inst_req_1); -- 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => array_obj_ref_1706_index_offset_req_1); -- 
    req_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => addr_of_1707_final_reg_req_1); -- 
    cr_4230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => ptr_deref_1711_load_0_req_1); -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => array_obj_ref_1729_index_offset_req_1); -- 
    req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => addr_of_1730_final_reg_req_1); -- 
    cr_4331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => ptr_deref_1733_store_0_req_1); -- 
    rr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1738_inst_req_0); -- 
    cr_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1738_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(98) & convTransposeA_CP_3758_elements(99) & convTransposeA_CP_3758_elements(100) & convTransposeA_CP_3758_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/$exit
      -- 
    ra_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => convTransposeA_CP_3758_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/$exit
      -- 
    ca_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => convTransposeA_CP_3758_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/$exit
      -- CP-element group 105: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/$exit
      -- CP-element group 105: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_req
      -- 
    phi_stmt_1822_req_4626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1822_req_4626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(105), ack => phi_stmt_1822_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(103) & convTransposeA_CP_3758_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Sample/$exit
      -- 
    ra_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_0, ack => convTransposeA_CP_3758_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/Update/ca
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1819_inst_ack_1, ack => convTransposeA_CP_3758_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- CP-element group 108: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1819/$exit
      -- CP-element group 108: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1816/$exit
      -- 
    phi_stmt_1816_req_4649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_4649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(108), ack => phi_stmt_1816_req_0); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(106) & convTransposeA_CP_3758_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/$exit
      -- CP-element group 109: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_req
      -- CP-element group 109: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1813_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/$exit
      -- 
    phi_stmt_1809_req_4657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1809_req_4657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(109), ack => phi_stmt_1809_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(76), ack => convTransposeA_CP_3758_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1491/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(105) & convTransposeA_CP_3758_elements(108) & convTransposeA_CP_3758_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/$exit
      -- 
    ra_4677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_0, ack => convTransposeA_CP_3758_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/$exit
      -- 
    ca_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_1, ack => convTransposeA_CP_3758_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_req
      -- CP-element group 113: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/$exit
      -- CP-element group 113: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/$exit
      -- 
    phi_stmt_1822_req_4683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1822_req_4683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(113), ack => phi_stmt_1822_req_1); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(111) & convTransposeA_CP_3758_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Sample/ra
      -- 
    ra_4700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_0, ack => convTransposeA_CP_3758_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/Update/$exit
      -- 
    ca_4705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_1, ack => convTransposeA_CP_3758_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/$exit
      -- CP-element group 116: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_req
      -- CP-element group 116: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1816/phi_stmt_1816_sources/type_cast_1821/$exit
      -- 
    phi_stmt_1816_req_4706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1816_req_4706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(116), ack => phi_stmt_1816_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(114) & convTransposeA_CP_3758_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Sample/ra
      -- 
    ra_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_0, ack => convTransposeA_CP_3758_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/Update/ca
      -- 
    ca_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_1, ack => convTransposeA_CP_3758_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/$exit
      -- CP-element group 119: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_req
      -- CP-element group 119: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1809/phi_stmt_1809_sources/type_cast_1815/$exit
      -- 
    phi_stmt_1809_req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1809_req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(119), ack => phi_stmt_1809_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(117) & convTransposeA_CP_3758_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1491/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(113) & convTransposeA_CP_3758_elements(116) & convTransposeA_CP_3758_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1491/merge_stmt_1808_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1491/merge_stmt_1808_PhiAck/$entry
      -- 
    convTransposeA_CP_3758_elements(121) <= OrReduce(convTransposeA_CP_3758_elements(110) & convTransposeA_CP_3758_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1491/merge_stmt_1808_PhiAck/phi_stmt_1809_ack
      -- 
    phi_stmt_1809_ack_4734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1809_ack_0, ack => convTransposeA_CP_3758_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1491/merge_stmt_1808_PhiAck/phi_stmt_1816_ack
      -- 
    phi_stmt_1816_ack_4735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1816_ack_0, ack => convTransposeA_CP_3758_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1491/merge_stmt_1808_PhiAck/phi_stmt_1822_ack
      -- 
    phi_stmt_1822_ack_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1822_ack_0, ack => convTransposeA_CP_3758_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1491/merge_stmt_1808_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(122) & convTransposeA_CP_3758_elements(123) & convTransposeA_CP_3758_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1728_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1728_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1705_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1705_scaled : std_logic_vector(13 downto 0);
    signal add41_1559 : std_logic_vector(15 downto 0);
    signal add54_1570 : std_logic_vector(15 downto 0);
    signal add73_1681 : std_logic_vector(63 downto 0);
    signal add75_1691 : std_logic_vector(63 downto 0);
    signal add86_1745 : std_logic_vector(31 downto 0);
    signal add93_1763 : std_logic_vector(15 downto 0);
    signal add_1543 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1639 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1706_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1706_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1706_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1706_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1706_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1706_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1708 : std_logic_vector(31 downto 0);
    signal arrayidx82_1731 : std_logic_vector(31 downto 0);
    signal call11_1512 : std_logic_vector(15 downto 0);
    signal call13_1515 : std_logic_vector(15 downto 0);
    signal call14_1518 : std_logic_vector(15 downto 0);
    signal call15_1521 : std_logic_vector(15 downto 0);
    signal call16_1534 : std_logic_vector(15 downto 0);
    signal call18_1546 : std_logic_vector(15 downto 0);
    signal call1_1497 : std_logic_vector(15 downto 0);
    signal call20_1549 : std_logic_vector(15 downto 0);
    signal call22_1552 : std_logic_vector(15 downto 0);
    signal call3_1500 : std_logic_vector(15 downto 0);
    signal call5_1503 : std_logic_vector(15 downto 0);
    signal call7_1506 : std_logic_vector(15 downto 0);
    signal call9_1509 : std_logic_vector(15 downto 0);
    signal call_1494 : std_logic_vector(15 downto 0);
    signal cmp101_1776 : std_logic_vector(0 downto 0);
    signal cmp112_1801 : std_logic_vector(0 downto 0);
    signal cmp_1750 : std_logic_vector(0 downto 0);
    signal conv107_1796 : std_logic_vector(31 downto 0);
    signal conv110_1591 : std_logic_vector(31 downto 0);
    signal conv17_1538 : std_logic_vector(31 downto 0);
    signal conv61_1663 : std_logic_vector(63 downto 0);
    signal conv64_1579 : std_logic_vector(63 downto 0);
    signal conv66_1667 : std_logic_vector(63 downto 0);
    signal conv69_1583 : std_logic_vector(63 downto 0);
    signal conv71_1671 : std_logic_vector(63 downto 0);
    signal conv85_1739 : std_logic_vector(31 downto 0);
    signal conv89_1587 : std_logic_vector(31 downto 0);
    signal conv_1525 : std_logic_vector(31 downto 0);
    signal idxprom81_1724 : std_logic_vector(63 downto 0);
    signal idxprom_1701 : std_logic_vector(63 downto 0);
    signal inc105_1780 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1785 : std_logic_vector(15 downto 0);
    signal inc_1771 : std_logic_vector(15 downto 0);
    signal indvar_1600 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1834 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1822 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1621 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1816 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1614 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1792 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1809 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1607 : std_logic_vector(15 downto 0);
    signal mul50_1654 : std_logic_vector(15 downto 0);
    signal mul72_1676 : std_logic_vector(63 downto 0);
    signal mul74_1686 : std_logic_vector(63 downto 0);
    signal mul_1644 : std_logic_vector(15 downto 0);
    signal ptr_deref_1711_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1711_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1711_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1711_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1711_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1733_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1733_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1531 : std_logic_vector(31 downto 0);
    signal shr111126_1597 : std_logic_vector(31 downto 0);
    signal shr80_1718 : std_logic_vector(63 downto 0);
    signal shr_1697 : std_logic_vector(31 downto 0);
    signal sub44_1649 : std_logic_vector(15 downto 0);
    signal sub57_1575 : std_logic_vector(15 downto 0);
    signal sub58_1659 : std_logic_vector(15 downto 0);
    signal sub_1564 : std_logic_vector(15 downto 0);
    signal tmp1_1634 : std_logic_vector(31 downto 0);
    signal tmp78_1712 : std_logic_vector(63 downto 0);
    signal type_cast_1529_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1557_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1595_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1606_wire : std_logic_vector(31 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1613_wire : std_logic_vector(15 downto 0);
    signal type_cast_1618_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1620_wire : std_logic_vector(15 downto 0);
    signal type_cast_1625_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1627_wire : std_logic_vector(15 downto 0);
    signal type_cast_1632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1695_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1722_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1743_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1761_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1769_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1789_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1813_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1815_wire : std_logic_vector(15 downto 0);
    signal type_cast_1819_wire : std_logic_vector(15 downto 0);
    signal type_cast_1821_wire : std_logic_vector(15 downto 0);
    signal type_cast_1825_wire : std_logic_vector(15 downto 0);
    signal type_cast_1827_wire : std_logic_vector(15 downto 0);
    signal type_cast_1832_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1840_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1706_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1706_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1706_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1706_resized_base_address <= "00000000000000";
    array_obj_ref_1729_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1729_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1729_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1729_resized_base_address <= "00000000000000";
    ptr_deref_1711_word_offset_0 <= "00000000000000";
    ptr_deref_1733_word_offset_0 <= "00000000000000";
    type_cast_1529_wire_constant <= "00000000000000000000000000010000";
    type_cast_1557_wire_constant <= "1111111111111111";
    type_cast_1568_wire_constant <= "1111111111111111";
    type_cast_1595_wire_constant <= "00000000000000000000000000000010";
    type_cast_1604_wire_constant <= "00000000000000000000000000000000";
    type_cast_1611_wire_constant <= "0000000000000000";
    type_cast_1618_wire_constant <= "0000000000000000";
    type_cast_1625_wire_constant <= "0000000000000000";
    type_cast_1632_wire_constant <= "00000000000000000000000000000100";
    type_cast_1695_wire_constant <= "00000000000000000000000000000010";
    type_cast_1716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1722_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1743_wire_constant <= "00000000000000000000000000000100";
    type_cast_1761_wire_constant <= "0000000000000100";
    type_cast_1769_wire_constant <= "0000000000000001";
    type_cast_1789_wire_constant <= "0000000000000000";
    type_cast_1813_wire_constant <= "0000000000000000";
    type_cast_1832_wire_constant <= "00000000000000000000000000000001";
    type_cast_1840_wire_constant <= "0000000000000001";
    phi_stmt_1600: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1604_wire_constant & type_cast_1606_wire;
      req <= phi_stmt_1600_req_0 & phi_stmt_1600_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1600",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1600_ack_0,
          idata => idata,
          odata => indvar_1600,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1600
    phi_stmt_1607: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1611_wire_constant & type_cast_1613_wire;
      req <= phi_stmt_1607_req_0 & phi_stmt_1607_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1607",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1607_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1607,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1607
    phi_stmt_1614: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1618_wire_constant & type_cast_1620_wire;
      req <= phi_stmt_1614_req_0 & phi_stmt_1614_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1614",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1614_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1614,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1614
    phi_stmt_1621: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1625_wire_constant & type_cast_1627_wire;
      req <= phi_stmt_1621_req_0 & phi_stmt_1621_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1621",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1621_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1621,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1621
    phi_stmt_1809: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1813_wire_constant & type_cast_1815_wire;
      req <= phi_stmt_1809_req_0 & phi_stmt_1809_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1809",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1809_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1809,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1809
    phi_stmt_1816: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1819_wire & type_cast_1821_wire;
      req <= phi_stmt_1816_req_0 & phi_stmt_1816_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1816",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1816_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1816,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1816
    phi_stmt_1822: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1825_wire & type_cast_1827_wire;
      req <= phi_stmt_1822_req_0 & phi_stmt_1822_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1822",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1822_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1822,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1822
    -- flow-through select operator MUX_1791_inst
    input_dim1x_x2_1792 <= type_cast_1789_wire_constant when (cmp101_1776(0) /=  '0') else inc_1771;
    addr_of_1707_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1707_final_reg_req_0;
      addr_of_1707_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1707_final_reg_req_1;
      addr_of_1707_final_reg_ack_1<= rack(0);
      addr_of_1707_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1707_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1706_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1730_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1730_final_reg_req_0;
      addr_of_1730_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1730_final_reg_req_1;
      addr_of_1730_final_reg_ack_1<= rack(0);
      addr_of_1730_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1730_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1729_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1524_inst_req_0;
      type_cast_1524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1524_inst_req_1;
      type_cast_1524_inst_ack_1<= rack(0);
      type_cast_1524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1524_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1521,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1525,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1537_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1537_inst_req_0;
      type_cast_1537_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1537_inst_req_1;
      type_cast_1537_inst_ack_1<= rack(0);
      type_cast_1537_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1537_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1534,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1578_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1578_inst_req_0;
      type_cast_1578_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1578_inst_req_1;
      type_cast_1578_inst_ack_1<= rack(0);
      type_cast_1578_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1578_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1552,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1579,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1582_inst_req_0;
      type_cast_1582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1582_inst_req_1;
      type_cast_1582_inst_ack_1<= rack(0);
      type_cast_1582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1549,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1586_inst_req_0;
      type_cast_1586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1586_inst_req_1;
      type_cast_1586_inst_ack_1<= rack(0);
      type_cast_1586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1587,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1590_inst_req_0;
      type_cast_1590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1590_inst_req_1;
      type_cast_1590_inst_ack_1<= rack(0);
      type_cast_1590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack(0);
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1809,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1613_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1620_inst_req_0;
      type_cast_1620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1620_inst_req_1;
      type_cast_1620_inst_ack_1<= rack(0);
      type_cast_1620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1816,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1620_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1627_inst_req_0;
      type_cast_1627_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1627_inst_req_1;
      type_cast_1627_inst_ack_1<= rack(0);
      type_cast_1627_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1627_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1627_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1662_inst_req_0;
      type_cast_1662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1662_inst_req_1;
      type_cast_1662_inst_ack_1<= rack(0);
      type_cast_1662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1662_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1663,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1666_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1666_inst_req_0;
      type_cast_1666_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1666_inst_req_1;
      type_cast_1666_inst_ack_1<= rack(0);
      type_cast_1666_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1666_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1667,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1670_inst_req_0;
      type_cast_1670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1670_inst_req_1;
      type_cast_1670_inst_ack_1<= rack(0);
      type_cast_1670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1700_inst_req_0;
      type_cast_1700_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1700_inst_req_1;
      type_cast_1700_inst_ack_1<= rack(0);
      type_cast_1700_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1700_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1697,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1701,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1738_inst_req_0;
      type_cast_1738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1738_inst_req_1;
      type_cast_1738_inst_ack_1<= rack(0);
      type_cast_1738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1739,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1779_inst_req_0;
      type_cast_1779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1779_inst_req_1;
      type_cast_1779_inst_ack_1<= rack(0);
      type_cast_1779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1795_inst_req_0;
      type_cast_1795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1795_inst_req_1;
      type_cast_1795_inst_ack_1<= rack(0);
      type_cast_1795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1785,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1815_inst_req_0;
      type_cast_1815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1815_inst_req_1;
      type_cast_1815_inst_ack_1<= rack(0);
      type_cast_1815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1763,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1815_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1819_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1819_inst_req_0;
      type_cast_1819_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1819_inst_req_1;
      type_cast_1819_inst_ack_1<= rack(0);
      type_cast_1819_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1819_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1819_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1821_inst_req_0;
      type_cast_1821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1821_inst_req_1;
      type_cast_1821_inst_ack_1<= rack(0);
      type_cast_1821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1821_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1785,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1825_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1827_inst_req_0;
      type_cast_1827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1827_inst_req_1;
      type_cast_1827_inst_ack_1<= rack(0);
      type_cast_1827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1827_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1706_index_1_rename
    process(R_idxprom_1705_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1705_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1705_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1706_index_1_resize
    process(idxprom_1701) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1701;
      ov := iv(13 downto 0);
      R_idxprom_1705_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1706_root_address_inst
    process(array_obj_ref_1706_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1706_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1706_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_index_1_rename
    process(R_idxprom81_1728_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1728_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1728_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_index_1_resize
    process(idxprom81_1724) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1724;
      ov := iv(13 downto 0);
      R_idxprom81_1728_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_root_address_inst
    process(array_obj_ref_1729_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1729_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1729_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1711_addr_0
    process(ptr_deref_1711_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1711_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1711_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1711_base_resize
    process(arrayidx77_1708) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1708;
      ov := iv(13 downto 0);
      ptr_deref_1711_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1711_gather_scatter
    process(ptr_deref_1711_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1711_data_0;
      ov(63 downto 0) := iv;
      tmp78_1712 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1711_root_address_inst
    process(ptr_deref_1711_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1711_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1711_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_addr_0
    process(ptr_deref_1733_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1733_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1733_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_base_resize
    process(arrayidx82_1731) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1731;
      ov := iv(13 downto 0);
      ptr_deref_1733_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_gather_scatter
    process(tmp78_1712) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1712;
      ov(63 downto 0) := iv;
      ptr_deref_1733_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_root_address_inst
    process(ptr_deref_1733_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1733_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1733_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1751_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1750;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1751_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1751_branch_req_0,
          ack0 => if_stmt_1751_branch_ack_0,
          ack1 => if_stmt_1751_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1802_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1801;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1802_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1802_branch_req_0,
          ack0 => if_stmt_1802_branch_ack_0,
          ack1 => if_stmt_1802_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1558_inst
    process(call7_1506) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1506, type_cast_1557_wire_constant, tmp_var);
      add41_1559 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1569_inst
    process(call9_1509) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1509, type_cast_1568_wire_constant, tmp_var);
      add54_1570 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1648_inst
    process(sub_1564, mul_1644) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1564, mul_1644, tmp_var);
      sub44_1649 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1658_inst
    process(sub57_1575, mul50_1654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1575, mul50_1654, tmp_var);
      sub58_1659 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1762_inst
    process(input_dim2x_x1_1607) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1607, type_cast_1761_wire_constant, tmp_var);
      add93_1763 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1770_inst
    process(input_dim1x_x1_1614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1614, type_cast_1769_wire_constant, tmp_var);
      inc_1771 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1784_inst
    process(inc105_1780, input_dim0x_x2_1621) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1780, input_dim0x_x2_1621, tmp_var);
      inc105x_xinput_dim0x_x2_1785 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1638_inst
    process(add_1543, tmp1_1634) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1543, tmp1_1634, tmp_var);
      add_src_0x_x0_1639 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1744_inst
    process(conv85_1739) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1739, type_cast_1743_wire_constant, tmp_var);
      add86_1745 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1833_inst
    process(indvar_1600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1600, type_cast_1832_wire_constant, tmp_var);
      indvarx_xnext_1834 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1680_inst
    process(mul72_1676, conv66_1667) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1676, conv66_1667, tmp_var);
      add73_1681 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1690_inst
    process(mul74_1686, conv61_1663) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1686, conv61_1663, tmp_var);
      add75_1691 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1723_inst
    process(shr80_1718) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1718, type_cast_1722_wire_constant, tmp_var);
      idxprom81_1724 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1775_inst
    process(inc_1771, call1_1497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1771, call1_1497, tmp_var);
      cmp101_1776 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1800_inst
    process(conv107_1796, shr111126_1597) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1796, shr111126_1597, tmp_var);
      cmp112_1801 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1596_inst
    process(conv110_1591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1591, type_cast_1595_wire_constant, tmp_var);
      shr111126_1597 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1696_inst
    process(add_src_0x_x0_1639) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1639, type_cast_1695_wire_constant, tmp_var);
      shr_1697 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1717_inst
    process(add75_1691) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1691, type_cast_1716_wire_constant, tmp_var);
      shr80_1718 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1643_inst
    process(input_dim0x_x2_1621, call13_1515) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1621, call13_1515, tmp_var);
      mul_1644 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1653_inst
    process(input_dim1x_x1_1614, call13_1515) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1614, call13_1515, tmp_var);
      mul50_1654 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1633_inst
    process(indvar_1600) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1600, type_cast_1632_wire_constant, tmp_var);
      tmp1_1634 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1675_inst
    process(conv71_1671, conv69_1583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1671, conv69_1583, tmp_var);
      mul72_1676 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1685_inst
    process(add73_1681, conv64_1579) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1681, conv64_1579, tmp_var);
      mul74_1686 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1542_inst
    process(shl_1531, conv17_1538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1531, conv17_1538, tmp_var);
      add_1543 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1530_inst
    process(conv_1525) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1525, type_cast_1529_wire_constant, tmp_var);
      shl_1531 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1563_inst
    process(add41_1559, call14_1518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1559, call14_1518, tmp_var);
      sub_1564 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1574_inst
    process(add54_1570, call14_1518) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1570, call14_1518, tmp_var);
      sub57_1575 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1749_inst
    process(add86_1745, conv89_1587) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1745, conv89_1587, tmp_var);
      cmp_1750 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1706_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1705_scaled;
      array_obj_ref_1706_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1706_index_offset_req_0;
      array_obj_ref_1706_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1706_index_offset_req_1;
      array_obj_ref_1706_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1729_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1728_scaled;
      array_obj_ref_1729_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1729_index_offset_req_0;
      array_obj_ref_1729_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1729_index_offset_req_1;
      array_obj_ref_1729_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1711_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1711_load_0_req_0;
      ptr_deref_1711_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1711_load_0_req_1;
      ptr_deref_1711_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1711_word_address_0;
      ptr_deref_1711_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1733_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1733_store_0_req_0;
      ptr_deref_1733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1733_store_0_req_1;
      ptr_deref_1733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1733_word_address_0;
      data_in <= ptr_deref_1733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1533_inst RPIPE_Block0_start_1545_inst RPIPE_Block0_start_1548_inst RPIPE_Block0_start_1551_inst RPIPE_Block0_start_1496_inst RPIPE_Block0_start_1499_inst RPIPE_Block0_start_1502_inst RPIPE_Block0_start_1505_inst RPIPE_Block0_start_1493_inst RPIPE_Block0_start_1508_inst RPIPE_Block0_start_1511_inst RPIPE_Block0_start_1520_inst RPIPE_Block0_start_1517_inst RPIPE_Block0_start_1514_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1533_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1545_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1548_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1551_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1496_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1499_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1502_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1505_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1493_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1508_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1511_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1520_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1517_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1514_inst_req_0;
      RPIPE_Block0_start_1533_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1545_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1548_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1551_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1496_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1499_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1502_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1505_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1493_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1508_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1511_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1520_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1517_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1514_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1533_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1545_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1548_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1551_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1496_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1499_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1502_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1505_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1493_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1508_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1511_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1520_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1517_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1514_inst_req_1;
      RPIPE_Block0_start_1533_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1545_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1548_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1551_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1496_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1499_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1502_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1505_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1493_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1508_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1511_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1520_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1517_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1514_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call16_1534 <= data_out(223 downto 208);
      call18_1546 <= data_out(207 downto 192);
      call20_1549 <= data_out(191 downto 176);
      call22_1552 <= data_out(175 downto 160);
      call1_1497 <= data_out(159 downto 144);
      call3_1500 <= data_out(143 downto 128);
      call5_1503 <= data_out(127 downto 112);
      call7_1506 <= data_out(111 downto 96);
      call_1494 <= data_out(95 downto 80);
      call9_1509 <= data_out(79 downto 64);
      call11_1512 <= data_out(63 downto 48);
      call15_1521 <= data_out(47 downto 32);
      call14_1518 <= data_out(31 downto 16);
      call13_1515 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1838_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1838_inst_req_0;
      WPIPE_Block0_done_1838_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1838_inst_req_1;
      WPIPE_Block0_done_1838_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1840_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4753_start: Boolean;
  signal convTransposeB_CP_4753_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1870_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1861_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_1 : boolean;
  signal type_cast_2182_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1889_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1889_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1861_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1864_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1864_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1849_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1849_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1901_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1904_inst_ack_1 : boolean;
  signal phi_stmt_2177_ack_0 : boolean;
  signal type_cast_1893_inst_ack_0 : boolean;
  signal type_cast_1893_inst_req_0 : boolean;
  signal phi_stmt_2183_ack_0 : boolean;
  signal phi_stmt_2170_ack_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_1 : boolean;
  signal type_cast_2182_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1901_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1901_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1858_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1861_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1861_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1901_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1870_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1889_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_1 : boolean;
  signal type_cast_1893_inst_req_1 : boolean;
  signal type_cast_1893_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1889_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1852_inst_req_1 : boolean;
  signal type_cast_2188_inst_req_1 : boolean;
  signal type_cast_2023_inst_ack_0 : boolean;
  signal type_cast_1952_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_1 : boolean;
  signal type_cast_1952_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_1 : boolean;
  signal type_cast_1952_inst_req_0 : boolean;
  signal type_cast_1952_inst_ack_0 : boolean;
  signal type_cast_1880_inst_ack_1 : boolean;
  signal phi_stmt_2183_req_1 : boolean;
  signal type_cast_1880_inst_req_1 : boolean;
  signal type_cast_1948_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_0 : boolean;
  signal type_cast_1948_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_0 : boolean;
  signal type_cast_1880_inst_ack_0 : boolean;
  signal type_cast_1944_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_0 : boolean;
  signal type_cast_1880_inst_req_0 : boolean;
  signal type_cast_1948_inst_req_0 : boolean;
  signal type_cast_1948_inst_ack_0 : boolean;
  signal type_cast_2023_inst_req_0 : boolean;
  signal type_cast_2188_inst_ack_1 : boolean;
  signal type_cast_1944_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_ack_1 : boolean;
  signal type_cast_1944_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_req_1 : boolean;
  signal type_cast_1944_inst_req_0 : boolean;
  signal type_cast_2023_inst_req_1 : boolean;
  signal type_cast_2023_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1904_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1904_inst_req_1 : boolean;
  signal type_cast_1940_inst_req_1 : boolean;
  signal type_cast_1940_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1849_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1904_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1864_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1849_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1864_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_0 : boolean;
  signal type_cast_1940_inst_req_0 : boolean;
  signal type_cast_1940_inst_ack_0 : boolean;
  signal type_cast_2027_inst_req_0 : boolean;
  signal type_cast_2027_inst_ack_0 : boolean;
  signal type_cast_2027_inst_req_1 : boolean;
  signal type_cast_2027_inst_ack_1 : boolean;
  signal type_cast_2188_inst_ack_0 : boolean;
  signal type_cast_2031_inst_req_0 : boolean;
  signal type_cast_2031_inst_ack_0 : boolean;
  signal type_cast_2031_inst_req_1 : boolean;
  signal type_cast_2031_inst_ack_1 : boolean;
  signal type_cast_2188_inst_req_0 : boolean;
  signal type_cast_2061_inst_req_0 : boolean;
  signal type_cast_2061_inst_ack_0 : boolean;
  signal type_cast_2061_inst_req_1 : boolean;
  signal type_cast_2061_inst_ack_1 : boolean;
  signal array_obj_ref_2067_index_offset_req_0 : boolean;
  signal array_obj_ref_2067_index_offset_ack_0 : boolean;
  signal array_obj_ref_2067_index_offset_req_1 : boolean;
  signal array_obj_ref_2067_index_offset_ack_1 : boolean;
  signal phi_stmt_2170_req_1 : boolean;
  signal addr_of_2068_final_reg_req_0 : boolean;
  signal addr_of_2068_final_reg_ack_0 : boolean;
  signal addr_of_2068_final_reg_req_1 : boolean;
  signal addr_of_2068_final_reg_ack_1 : boolean;
  signal ptr_deref_2072_load_0_req_0 : boolean;
  signal ptr_deref_2072_load_0_ack_0 : boolean;
  signal type_cast_2182_inst_ack_0 : boolean;
  signal ptr_deref_2072_load_0_req_1 : boolean;
  signal ptr_deref_2072_load_0_ack_1 : boolean;
  signal phi_stmt_2170_req_0 : boolean;
  signal type_cast_2173_inst_ack_1 : boolean;
  signal type_cast_2173_inst_req_1 : boolean;
  signal array_obj_ref_2090_index_offset_req_0 : boolean;
  signal array_obj_ref_2090_index_offset_ack_0 : boolean;
  signal array_obj_ref_2090_index_offset_req_1 : boolean;
  signal array_obj_ref_2090_index_offset_ack_1 : boolean;
  signal type_cast_2173_inst_ack_0 : boolean;
  signal addr_of_2091_final_reg_req_0 : boolean;
  signal addr_of_2091_final_reg_ack_0 : boolean;
  signal addr_of_2091_final_reg_req_1 : boolean;
  signal addr_of_2091_final_reg_ack_1 : boolean;
  signal type_cast_2173_inst_req_0 : boolean;
  signal phi_stmt_2183_req_0 : boolean;
  signal ptr_deref_2094_store_0_req_0 : boolean;
  signal ptr_deref_2094_store_0_ack_0 : boolean;
  signal type_cast_2182_inst_req_0 : boolean;
  signal type_cast_2186_inst_ack_1 : boolean;
  signal ptr_deref_2094_store_0_req_1 : boolean;
  signal ptr_deref_2094_store_0_ack_1 : boolean;
  signal type_cast_2099_inst_req_0 : boolean;
  signal type_cast_2099_inst_ack_0 : boolean;
  signal type_cast_2099_inst_req_1 : boolean;
  signal type_cast_2099_inst_ack_1 : boolean;
  signal if_stmt_2112_branch_req_0 : boolean;
  signal if_stmt_2112_branch_ack_1 : boolean;
  signal if_stmt_2112_branch_ack_0 : boolean;
  signal type_cast_2186_inst_req_1 : boolean;
  signal type_cast_2140_inst_req_0 : boolean;
  signal type_cast_2140_inst_ack_0 : boolean;
  signal type_cast_2140_inst_req_1 : boolean;
  signal type_cast_2140_inst_ack_1 : boolean;
  signal type_cast_2156_inst_req_0 : boolean;
  signal type_cast_2156_inst_ack_0 : boolean;
  signal type_cast_2156_inst_req_1 : boolean;
  signal type_cast_2156_inst_ack_1 : boolean;
  signal if_stmt_2163_branch_req_0 : boolean;
  signal if_stmt_2163_branch_ack_1 : boolean;
  signal if_stmt_2163_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2199_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2199_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2199_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2199_inst_ack_1 : boolean;
  signal type_cast_2186_inst_ack_0 : boolean;
  signal type_cast_1986_inst_req_0 : boolean;
  signal type_cast_1986_inst_ack_0 : boolean;
  signal type_cast_1986_inst_req_1 : boolean;
  signal type_cast_1986_inst_ack_1 : boolean;
  signal phi_stmt_1983_req_0 : boolean;
  signal phi_stmt_1976_req_0 : boolean;
  signal phi_stmt_1969_req_0 : boolean;
  signal phi_stmt_1962_req_1 : boolean;
  signal type_cast_2186_inst_req_0 : boolean;
  signal type_cast_1988_inst_req_0 : boolean;
  signal type_cast_1988_inst_ack_0 : boolean;
  signal phi_stmt_2177_req_0 : boolean;
  signal type_cast_1988_inst_req_1 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal type_cast_1988_inst_ack_1 : boolean;
  signal phi_stmt_1983_req_1 : boolean;
  signal type_cast_1982_inst_req_0 : boolean;
  signal type_cast_1982_inst_ack_0 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal type_cast_1982_inst_req_1 : boolean;
  signal type_cast_1982_inst_ack_1 : boolean;
  signal phi_stmt_1976_req_1 : boolean;
  signal type_cast_1975_inst_req_0 : boolean;
  signal type_cast_1975_inst_ack_0 : boolean;
  signal type_cast_1975_inst_req_1 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal type_cast_1975_inst_ack_1 : boolean;
  signal phi_stmt_1969_req_1 : boolean;
  signal type_cast_1965_inst_req_0 : boolean;
  signal type_cast_1965_inst_ack_0 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal type_cast_1965_inst_req_1 : boolean;
  signal type_cast_1965_inst_ack_1 : boolean;
  signal phi_stmt_1962_req_0 : boolean;
  signal phi_stmt_1962_ack_0 : boolean;
  signal phi_stmt_1969_ack_0 : boolean;
  signal phi_stmt_1976_ack_0 : boolean;
  signal phi_stmt_1983_ack_0 : boolean;
  signal phi_stmt_2177_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4753_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4753: Block -- control-path 
    signal convTransposeB_CP_4753_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4753_elements(0) <= convTransposeB_CP_4753_start;
    convTransposeB_CP_4753_symbol <= convTransposeB_CP_4753_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1847/branch_block_stmt_1847__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908__entry__
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1847/$entry
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/$entry
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Update/cr
      -- 
    rr_4801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => RPIPE_Block1_start_1849_inst_req_0); -- 
    cr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => type_cast_1893_inst_req_1); -- 
    cr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => type_cast_1880_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1847/assign_stmt_2195__exit__
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1847/assign_stmt_2195__entry__
      -- CP-element group 1: 	 branch_block_stmt_1847/merge_stmt_2169__exit__
      -- CP-element group 1: 	 branch_block_stmt_1847/assign_stmt_2195/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/assign_stmt_2195/$exit
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Update/cr
      -- 
    rr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1988_inst_req_0); -- 
    cr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1988_inst_req_1); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1982_inst_req_0); -- 
    cr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1982_inst_req_1); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1975_inst_req_0); -- 
    cr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1975_inst_req_1); -- 
    rr_5571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1965_inst_req_0); -- 
    cr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1965_inst_req_1); -- 
    convTransposeB_CP_4753_elements(1) <= convTransposeB_CP_4753_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Update/cr
      -- 
    ra_4802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1849_inst_ack_0, ack => convTransposeB_CP_4753_elements(2)); -- 
    cr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(2), ack => RPIPE_Block1_start_1849_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1849_Update/ca
      -- 
    ca_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1849_inst_ack_1, ack => convTransposeB_CP_4753_elements(3)); -- 
    rr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(3), ack => RPIPE_Block1_start_1852_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_sample_completed_
      -- 
    ra_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1852_inst_ack_0, ack => convTransposeB_CP_4753_elements(4)); -- 
    cr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(4), ack => RPIPE_Block1_start_1852_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1852_Update/$exit
      -- 
    ca_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1852_inst_ack_1, ack => convTransposeB_CP_4753_elements(5)); -- 
    rr_4829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(5), ack => RPIPE_Block1_start_1855_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_sample_completed_
      -- 
    ra_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_0, ack => convTransposeB_CP_4753_elements(6)); -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(6), ack => RPIPE_Block1_start_1855_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1855_update_completed_
      -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_1, ack => convTransposeB_CP_4753_elements(7)); -- 
    rr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(7), ack => RPIPE_Block1_start_1858_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Update/cr
      -- 
    ra_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1858_inst_ack_0, ack => convTransposeB_CP_4753_elements(8)); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(8), ack => RPIPE_Block1_start_1858_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1858_Update/$exit
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1858_inst_ack_1, ack => convTransposeB_CP_4753_elements(9)); -- 
    rr_4857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(9), ack => RPIPE_Block1_start_1861_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_sample_completed_
      -- 
    ra_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1861_inst_ack_0, ack => convTransposeB_CP_4753_elements(10)); -- 
    cr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(10), ack => RPIPE_Block1_start_1861_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1861_Update/ca
      -- 
    ca_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1861_inst_ack_1, ack => convTransposeB_CP_4753_elements(11)); -- 
    rr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(11), ack => RPIPE_Block1_start_1864_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Update/cr
      -- 
    ra_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1864_inst_ack_0, ack => convTransposeB_CP_4753_elements(12)); -- 
    cr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(12), ack => RPIPE_Block1_start_1864_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1864_Update/ca
      -- 
    ca_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1864_inst_ack_1, ack => convTransposeB_CP_4753_elements(13)); -- 
    rr_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(13), ack => RPIPE_Block1_start_1867_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_update_start_
      -- 
    ra_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_0, ack => convTransposeB_CP_4753_elements(14)); -- 
    cr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(14), ack => RPIPE_Block1_start_1867_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1867_update_completed_
      -- 
    ca_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_1, ack => convTransposeB_CP_4753_elements(15)); -- 
    rr_4899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(15), ack => RPIPE_Block1_start_1870_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_sample_completed_
      -- 
    ra_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_0, ack => convTransposeB_CP_4753_elements(16)); -- 
    cr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(16), ack => RPIPE_Block1_start_1870_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1870_Update/$exit
      -- 
    ca_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_1, ack => convTransposeB_CP_4753_elements(17)); -- 
    rr_4913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(17), ack => RPIPE_Block1_start_1873_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_sample_completed_
      -- 
    ra_4914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_0, ack => convTransposeB_CP_4753_elements(18)); -- 
    cr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(18), ack => RPIPE_Block1_start_1873_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1873_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Sample/$entry
      -- 
    ca_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_1, ack => convTransposeB_CP_4753_elements(19)); -- 
    rr_4927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(19), ack => RPIPE_Block1_start_1876_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Sample/$exit
      -- 
    ra_4928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_0, ack => convTransposeB_CP_4753_elements(20)); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(20), ack => RPIPE_Block1_start_1876_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1876_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Sample/$entry
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_1, ack => convTransposeB_CP_4753_elements(21)); -- 
    rr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(21), ack => type_cast_1880_inst_req_0); -- 
    rr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(21), ack => RPIPE_Block1_start_1889_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Sample/$exit
      -- 
    ra_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1880_inst_ack_0, ack => convTransposeB_CP_4753_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1880_update_completed_
      -- 
    ca_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1880_inst_ack_1, ack => convTransposeB_CP_4753_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_sample_completed_
      -- 
    ra_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1889_inst_ack_0, ack => convTransposeB_CP_4753_elements(24)); -- 
    cr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(24), ack => RPIPE_Block1_start_1889_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1889_update_completed_
      -- 
    ca_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1889_inst_ack_1, ack => convTransposeB_CP_4753_elements(25)); -- 
    rr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(25), ack => type_cast_1893_inst_req_0); -- 
    rr_4983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(25), ack => RPIPE_Block1_start_1901_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Sample/$exit
      -- 
    ra_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1893_inst_ack_0, ack => convTransposeB_CP_4753_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/type_cast_1893_Update/ca
      -- 
    ca_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1893_inst_ack_1, ack => convTransposeB_CP_4753_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Sample/$exit
      -- 
    ra_4984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1901_inst_ack_0, ack => convTransposeB_CP_4753_elements(28)); -- 
    cr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(28), ack => RPIPE_Block1_start_1901_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1901_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Sample/rr
      -- 
    ca_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1901_inst_ack_1, ack => convTransposeB_CP_4753_elements(29)); -- 
    rr_4997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(29), ack => RPIPE_Block1_start_1904_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Update/$entry
      -- 
    ra_4998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1904_inst_ack_0, ack => convTransposeB_CP_4753_elements(30)); -- 
    cr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(30), ack => RPIPE_Block1_start_1904_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1904_Update/$exit
      -- 
    ca_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1904_inst_ack_1, ack => convTransposeB_CP_4753_elements(31)); -- 
    rr_5011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(31), ack => RPIPE_Block1_start_1907_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Sample/ra
      -- 
    ra_5012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_0, ack => convTransposeB_CP_4753_elements(32)); -- 
    cr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(32), ack => RPIPE_Block1_start_1907_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/RPIPE_Block1_start_1907_Update/$exit
      -- 
    ca_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_1, ack => convTransposeB_CP_4753_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908__exit__
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1850_to_assign_stmt_1908/$exit
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959__entry__
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_sample_start_
      -- 
    cr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1952_inst_req_1); -- 
    rr_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1952_inst_req_0); -- 
    cr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1948_inst_req_1); -- 
    rr_5056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1948_inst_req_0); -- 
    cr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1944_inst_req_1); -- 
    rr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1944_inst_req_0); -- 
    cr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1940_inst_req_1); -- 
    rr_5028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1940_inst_req_0); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(23) & convTransposeB_CP_4753_elements(27) & convTransposeB_CP_4753_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_sample_completed_
      -- 
    ra_5029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1940_inst_ack_0, ack => convTransposeB_CP_4753_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1940_Update/$exit
      -- 
    ca_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1940_inst_ack_1, ack => convTransposeB_CP_4753_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_sample_completed_
      -- 
    ra_5043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_0, ack => convTransposeB_CP_4753_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1944_Update/$exit
      -- 
    ca_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_1, ack => convTransposeB_CP_4753_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_sample_completed_
      -- 
    ra_5057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1948_inst_ack_0, ack => convTransposeB_CP_4753_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1948_update_completed_
      -- 
    ca_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1948_inst_ack_1, ack => convTransposeB_CP_4753_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_sample_completed_
      -- 
    ra_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1952_inst_ack_0, ack => convTransposeB_CP_4753_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/type_cast_1952_update_completed_
      -- 
    ca_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1952_inst_ack_1, ack => convTransposeB_CP_4753_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959__exit__
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1847/assign_stmt_1915_to_assign_stmt_1959/$exit
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/$entry
      -- CP-element group 43: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/$entry
      -- 
    rr_5452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(43), ack => type_cast_1986_inst_req_0); -- 
    cr_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(43), ack => type_cast_1986_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(36) & convTransposeB_CP_4753_elements(38) & convTransposeB_CP_4753_elements(40) & convTransposeB_CP_4753_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Sample/$exit
      -- 
    ra_5088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_0, ack => convTransposeB_CP_4753_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Update/ca
      -- 
    ca_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_1, ack => convTransposeB_CP_4753_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Sample/ra
      -- 
    ra_5102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_0, ack => convTransposeB_CP_4753_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Update/ca
      -- 
    ca_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2027_inst_ack_1, ack => convTransposeB_CP_4753_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Sample/ra
      -- 
    ra_5116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_0, ack => convTransposeB_CP_4753_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Update/ca
      -- 
    ca_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2031_inst_ack_1, ack => convTransposeB_CP_4753_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Sample/ra
      -- 
    ra_5130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_0, ack => convTransposeB_CP_4753_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Sample/req
      -- 
    ca_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2061_inst_ack_1, ack => convTransposeB_CP_4753_elements(51)); -- 
    req_5160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(51), ack => array_obj_ref_2067_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Sample/ack
      -- 
    ack_5161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2067_index_offset_ack_0, ack => convTransposeB_CP_4753_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_request/req
      -- 
    ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2067_index_offset_ack_1, ack => convTransposeB_CP_4753_elements(53)); -- 
    req_5175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(53), ack => addr_of_2068_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_request/ack
      -- 
    ack_5176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2068_final_reg_ack_0, ack => convTransposeB_CP_4753_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/word_0/rr
      -- 
    ack_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2068_final_reg_ack_1, ack => convTransposeB_CP_4753_elements(55)); -- 
    rr_5214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(55), ack => ptr_deref_2072_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Sample/word_access_start/word_0/ra
      -- 
    ra_5215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2072_load_0_ack_0, ack => convTransposeB_CP_4753_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/ptr_deref_2072_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/ptr_deref_2072_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/ptr_deref_2072_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/ptr_deref_2072_Merge/merge_ack
      -- 
    ca_5226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2072_load_0_ack_1, ack => convTransposeB_CP_4753_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Sample/req
      -- 
    req_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(58), ack => array_obj_ref_2090_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(45) & convTransposeB_CP_4753_elements(47) & convTransposeB_CP_4753_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Sample/ack
      -- 
    ack_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2090_index_offset_ack_0, ack => convTransposeB_CP_4753_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_request/req
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2090_index_offset_ack_1, ack => convTransposeB_CP_4753_elements(60)); -- 
    req_5271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(60), ack => addr_of_2091_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_request/ack
      -- 
    ack_5272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2091_final_reg_ack_0, ack => convTransposeB_CP_4753_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_word_addrgen/root_register_ack
      -- 
    ack_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2091_final_reg_ack_1, ack => convTransposeB_CP_4753_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/ptr_deref_2094_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/ptr_deref_2094_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/ptr_deref_2094_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/ptr_deref_2094_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/word_0/rr
      -- 
    rr_5315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(63), ack => ptr_deref_2094_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(57) & convTransposeB_CP_4753_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Sample/word_access_start/word_0/ra
      -- 
    ra_5316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2094_store_0_ack_0, ack => convTransposeB_CP_4753_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/word_0/ca
      -- 
    ca_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2094_store_0_ack_1, ack => convTransposeB_CP_4753_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Sample/ra
      -- 
    ra_5336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2099_inst_ack_0, ack => convTransposeB_CP_4753_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Update/ca
      -- 
    ca_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2099_inst_ack_1, ack => convTransposeB_CP_4753_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111__exit__
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112__entry__
      -- CP-element group 68: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/$exit
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1847/R_cmp_2113_place
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1847/if_stmt_2112_else_link/$entry
      -- 
    branch_req_5349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(68), ack => if_stmt_2112_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(52) & convTransposeB_CP_4753_elements(59) & convTransposeB_CP_4753_elements(65) & convTransposeB_CP_4753_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/assign_stmt_2124__exit__
      -- CP-element group 69: 	 branch_block_stmt_1847/merge_stmt_2118__exit__
      -- CP-element group 69: 	 branch_block_stmt_1847/assign_stmt_2124__entry__
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/if_stmt_2112_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1847/if_stmt_2112_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1847/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1847/assign_stmt_2124/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/assign_stmt_2124/$exit
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1847/merge_stmt_2118_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1847/merge_stmt_2118_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1847/merge_stmt_2118_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1847/merge_stmt_2118_PhiAck/dummy
      -- 
    if_choice_transition_5354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_1, ack => convTransposeB_CP_4753_elements(69)); -- 
    cr_5737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2188_inst_req_1); -- 
    rr_5732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2188_inst_req_0); -- 
    cr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2173_inst_req_1); -- 
    rr_5709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2173_inst_req_0); -- 
    cr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2180_inst_req_1); -- 
    rr_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2180_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1847/merge_stmt_2126__exit__
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162__entry__
      -- CP-element group 70: 	 branch_block_stmt_1847/if_stmt_2112_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1847/if_stmt_2112_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1847/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/$entry
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1847/merge_stmt_2126_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1847/merge_stmt_2126_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1847/merge_stmt_2126_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1847/merge_stmt_2126_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1847/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1847/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- 
    else_choice_transition_5358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2112_branch_ack_0, ack => convTransposeB_CP_4753_elements(70)); -- 
    rr_5374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2140_inst_req_0); -- 
    cr_5379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2140_inst_req_1); -- 
    cr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2156_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Sample/ra
      -- 
    ra_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_0, ack => convTransposeB_CP_4753_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2140_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Sample/rr
      -- 
    ca_5380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_1, ack => convTransposeB_CP_4753_elements(72)); -- 
    rr_5388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(72), ack => type_cast_2156_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Sample/ra
      -- 
    ra_5389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2156_inst_ack_0, ack => convTransposeB_CP_4753_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162__exit__
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163__entry__
      -- CP-element group 74: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/$exit
      -- CP-element group 74: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1847/assign_stmt_2132_to_assign_stmt_2162/type_cast_2156_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1847/R_cmp117_2164_place
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1847/if_stmt_2163_else_link/$entry
      -- 
    ca_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2156_inst_ack_1, ack => convTransposeB_CP_4753_elements(74)); -- 
    branch_req_5402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(74), ack => if_stmt_2163_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1847/merge_stmt_2197__exit__
      -- CP-element group 75: 	 branch_block_stmt_1847/merge_stmt_2197_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1847/merge_stmt_2197_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1847/assign_stmt_2202__entry__
      -- CP-element group 75: 	 branch_block_stmt_1847/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1847/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1847/merge_stmt_2197_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1847/merge_stmt_2197_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1847/if_stmt_2163_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1847/if_stmt_2163_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1847/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1847/assign_stmt_2202/$entry
      -- CP-element group 75: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Sample/req
      -- 
    if_choice_transition_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2163_branch_ack_1, ack => convTransposeB_CP_4753_elements(75)); -- 
    req_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(75), ack => WPIPE_Block1_done_2199_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/if_stmt_2163_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/if_stmt_2163_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/$entry
      -- 
    else_choice_transition_5411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2163_branch_ack_0, ack => convTransposeB_CP_4753_elements(76)); -- 
    cr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2182_inst_req_1); -- 
    rr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2182_inst_req_0); -- 
    cr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2186_inst_req_1); -- 
    rr_5660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2186_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Update/req
      -- 
    ack_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2199_inst_ack_0, ack => convTransposeB_CP_4753_elements(77)); -- 
    req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(77), ack => WPIPE_Block1_done_2199_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1847/branch_block_stmt_1847__exit__
      -- CP-element group 78: 	 branch_block_stmt_1847/merge_stmt_2204_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1847/$exit
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1847/assign_stmt_2202__exit__
      -- CP-element group 78: 	 branch_block_stmt_1847/return__
      -- CP-element group 78: 	 branch_block_stmt_1847/merge_stmt_2204__exit__
      -- CP-element group 78: 	 branch_block_stmt_1847/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1847/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1847/merge_stmt_2204_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1847/assign_stmt_2202/$exit
      -- CP-element group 78: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1847/assign_stmt_2202/WPIPE_Block1_done_2199_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1847/merge_stmt_2204_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1847/merge_stmt_2204_PhiAck/$exit
      -- 
    ack_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2199_inst_ack_1, ack => convTransposeB_CP_4753_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Sample/ra
      -- 
    ra_5453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_0, ack => convTransposeB_CP_4753_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/Update/ca
      -- 
    ca_5458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1986_inst_ack_1, ack => convTransposeB_CP_4753_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/$exit
      -- CP-element group 81: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/$exit
      -- CP-element group 81: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1986/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_req
      -- 
    phi_stmt_1983_req_5459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_req_5459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(81), ack => phi_stmt_1983_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(79) & convTransposeB_CP_4753_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/$exit
      -- CP-element group 82: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1980_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_req
      -- 
    phi_stmt_1976_req_5467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1976_req_5467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(82), ack => phi_stmt_1976_req_0); -- 
    -- Element group convTransposeB_CP_4753_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/$exit
      -- CP-element group 83: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1973_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_req
      -- 
    phi_stmt_1969_req_5475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_req_5475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(83), ack => phi_stmt_1969_req_0); -- 
    -- Element group convTransposeB_CP_4753_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/$exit
      -- CP-element group 84: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1968_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_req
      -- 
    phi_stmt_1962_req_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1962_req_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(84), ack => phi_stmt_1962_req_1); -- 
    -- Element group convTransposeB_CP_4753_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1847/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(81) & convTransposeB_CP_4753_elements(82) & convTransposeB_CP_4753_elements(83) & convTransposeB_CP_4753_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Sample/ra
      -- 
    ra_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_0, ack => convTransposeB_CP_4753_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/Update/ca
      -- 
    ca_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1988_inst_ack_1, ack => convTransposeB_CP_4753_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/$exit
      -- CP-element group 88: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/$exit
      -- CP-element group 88: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_sources/type_cast_1988/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1983/phi_stmt_1983_req
      -- 
    phi_stmt_1983_req_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1983_req_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(88), ack => phi_stmt_1983_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(86) & convTransposeB_CP_4753_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Sample/ra
      -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1982_inst_ack_0, ack => convTransposeB_CP_4753_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/Update/ca
      -- 
    ca_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1982_inst_ack_1, ack => convTransposeB_CP_4753_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/$exit
      -- CP-element group 91: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/$exit
      -- CP-element group 91: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_sources/type_cast_1982/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1976/phi_stmt_1976_req
      -- 
    phi_stmt_1976_req_5532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1976_req_5532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(91), ack => phi_stmt_1976_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(89) & convTransposeB_CP_4753_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Sample/ra
      -- 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_0, ack => convTransposeB_CP_4753_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/Update/ca
      -- 
    ca_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_1, ack => convTransposeB_CP_4753_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/$exit
      -- CP-element group 94: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/$exit
      -- CP-element group 94: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_sources/type_cast_1975/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1969/phi_stmt_1969_req
      -- 
    phi_stmt_1969_req_5555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1969_req_5555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(94), ack => phi_stmt_1969_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(92) & convTransposeB_CP_4753_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Sample/ra
      -- 
    ra_5572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1965_inst_ack_0, ack => convTransposeB_CP_4753_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/Update/ca
      -- 
    ca_5577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1965_inst_ack_1, ack => convTransposeB_CP_4753_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/$exit
      -- CP-element group 97: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/$exit
      -- CP-element group 97: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_sources/type_cast_1965/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1962/phi_stmt_1962_req
      -- 
    phi_stmt_1962_req_5578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1962_req_5578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(97), ack => phi_stmt_1962_req_0); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(95) & convTransposeB_CP_4753_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1847/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(88) & convTransposeB_CP_4753_elements(91) & convTransposeB_CP_4753_elements(94) & convTransposeB_CP_4753_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1847/merge_stmt_1961_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/$entry
      -- 
    convTransposeB_CP_4753_elements(99) <= OrReduce(convTransposeB_CP_4753_elements(85) & convTransposeB_CP_4753_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/phi_stmt_1962_ack
      -- 
    phi_stmt_1962_ack_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1962_ack_0, ack => convTransposeB_CP_4753_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/phi_stmt_1969_ack
      -- 
    phi_stmt_1969_ack_5584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1969_ack_0, ack => convTransposeB_CP_4753_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/phi_stmt_1976_ack
      -- 
    phi_stmt_1976_ack_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1976_ack_0, ack => convTransposeB_CP_4753_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/phi_stmt_1983_ack
      -- 
    phi_stmt_1983_ack_5586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1983_ack_0, ack => convTransposeB_CP_4753_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1847/merge_stmt_1961__exit__
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111__entry__
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2023_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2027_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2031_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2061_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2067_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2068_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2072_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/array_obj_ref_2090_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/addr_of_2091_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/ptr_deref_2094_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1847/assign_stmt_1995_to_assign_stmt_2111/type_cast_2099_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1847/merge_stmt_1961_PhiAck/$exit
      -- 
    rr_5087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2023_inst_req_0); -- 
    cr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2023_inst_req_1); -- 
    rr_5101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2027_inst_req_0); -- 
    cr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2027_inst_req_1); -- 
    rr_5115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2031_inst_req_0); -- 
    cr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2031_inst_req_1); -- 
    rr_5129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2061_inst_req_0); -- 
    cr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2061_inst_req_1); -- 
    req_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => array_obj_ref_2067_index_offset_req_1); -- 
    req_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => addr_of_2068_final_reg_req_1); -- 
    cr_5225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => ptr_deref_2072_load_0_req_1); -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => array_obj_ref_2090_index_offset_req_1); -- 
    req_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => addr_of_2091_final_reg_req_1); -- 
    cr_5326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => ptr_deref_2094_store_0_req_1); -- 
    rr_5335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2099_inst_req_0); -- 
    cr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2099_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(100) & convTransposeB_CP_4753_elements(101) & convTransposeB_CP_4753_elements(102) & convTransposeB_CP_4753_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Sample/$exit
      -- 
    ra_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_0, ack => convTransposeB_CP_4753_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/Update/$exit
      -- 
    ca_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_1, ack => convTransposeB_CP_4753_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2182/$exit
      -- CP-element group 107: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/$exit
      -- CP-element group 107: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_req
      -- 
    phi_stmt_2177_req_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2177_req_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(107), ack => phi_stmt_2177_req_1); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(105) & convTransposeB_CP_4753_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_req
      -- CP-element group 108: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2176_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2170/$exit
      -- 
    phi_stmt_2170_req_5644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2170_req_5644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(108), ack => phi_stmt_2170_req_1); -- 
    -- Element group convTransposeB_CP_4753_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(76), ack => convTransposeB_CP_4753_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/$exit
      -- 
    ra_5661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_0, ack => convTransposeB_CP_4753_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/ca
      -- CP-element group 110: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/$exit
      -- 
    ca_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_1, ack => convTransposeB_CP_4753_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/$exit
      -- CP-element group 111: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/$exit
      -- CP-element group 111: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_req
      -- CP-element group 111: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/$exit
      -- 
    phi_stmt_2183_req_5667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2183_req_5667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(111), ack => phi_stmt_2183_req_0); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(109) & convTransposeB_CP_4753_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1847/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(107) & convTransposeB_CP_4753_elements(108) & convTransposeB_CP_4753_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Sample/$exit
      -- 
    ra_5687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => convTransposeB_CP_4753_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/Update/$exit
      -- 
    ca_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => convTransposeB_CP_4753_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/$exit
      -- CP-element group 115: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/$exit
      -- CP-element group 115: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_req
      -- CP-element group 115: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2177/phi_stmt_2177_sources/type_cast_2180/SplitProtocol/$exit
      -- 
    phi_stmt_2177_req_5693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2177_req_5693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(115), ack => phi_stmt_2177_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(113) & convTransposeB_CP_4753_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Sample/$exit
      -- 
    ra_5710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2173_inst_ack_0, ack => convTransposeB_CP_4753_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/Update/$exit
      -- 
    ca_5715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2173_inst_ack_1, ack => convTransposeB_CP_4753_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_req
      -- CP-element group 118: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/type_cast_2173/$exit
      -- CP-element group 118: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/phi_stmt_2170_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2170/$exit
      -- 
    phi_stmt_2170_req_5716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2170_req_5716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(118), ack => phi_stmt_2170_req_0); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(116) & convTransposeB_CP_4753_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/$exit
      -- 
    ra_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_0, ack => convTransposeB_CP_4753_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/$exit
      -- 
    ca_5738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_1, ack => convTransposeB_CP_4753_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_req
      -- CP-element group 121: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/$exit
      -- CP-element group 121: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/$exit
      -- 
    phi_stmt_2183_req_5739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2183_req_5739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(121), ack => phi_stmt_2183_req_1); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(119) & convTransposeB_CP_4753_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1847/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(115) & convTransposeB_CP_4753_elements(118) & convTransposeB_CP_4753_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1847/merge_stmt_2169_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_1847/merge_stmt_2169_PhiReqMerge
      -- 
    convTransposeB_CP_4753_elements(123) <= OrReduce(convTransposeB_CP_4753_elements(112) & convTransposeB_CP_4753_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1847/merge_stmt_2169_PhiAck/phi_stmt_2170_ack
      -- 
    phi_stmt_2170_ack_5744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2170_ack_0, ack => convTransposeB_CP_4753_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1847/merge_stmt_2169_PhiAck/phi_stmt_2177_ack
      -- 
    phi_stmt_2177_ack_5745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2177_ack_0, ack => convTransposeB_CP_4753_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1847/merge_stmt_2169_PhiAck/phi_stmt_2183_ack
      -- 
    phi_stmt_2183_ack_5746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2183_ack_0, ack => convTransposeB_CP_4753_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1847/merge_stmt_2169_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(124) & convTransposeB_CP_4753_elements(125) & convTransposeB_CP_4753_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2089_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2089_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2066_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2066_scaled : std_logic_vector(13 downto 0);
    signal add45_1921 : std_logic_vector(15 downto 0);
    signal add58_1932 : std_logic_vector(15 downto 0);
    signal add77_2042 : std_logic_vector(63 downto 0);
    signal add79_2052 : std_logic_vector(63 downto 0);
    signal add91_2106 : std_logic_vector(31 downto 0);
    signal add98_2124 : std_logic_vector(15 downto 0);
    signal add_1899 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2000 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2067_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2067_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2090_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2069 : std_logic_vector(31 downto 0);
    signal arrayidx87_2092 : std_logic_vector(31 downto 0);
    signal call11_1868 : std_logic_vector(15 downto 0);
    signal call13_1871 : std_logic_vector(15 downto 0);
    signal call14_1874 : std_logic_vector(15 downto 0);
    signal call15_1877 : std_logic_vector(15 downto 0);
    signal call16_1890 : std_logic_vector(15 downto 0);
    signal call18_1902 : std_logic_vector(15 downto 0);
    signal call1_1853 : std_logic_vector(15 downto 0);
    signal call20_1905 : std_logic_vector(15 downto 0);
    signal call22_1908 : std_logic_vector(15 downto 0);
    signal call3_1856 : std_logic_vector(15 downto 0);
    signal call5_1859 : std_logic_vector(15 downto 0);
    signal call7_1862 : std_logic_vector(15 downto 0);
    signal call9_1865 : std_logic_vector(15 downto 0);
    signal call_1850 : std_logic_vector(15 downto 0);
    signal cmp106_2137 : std_logic_vector(0 downto 0);
    signal cmp117_2162 : std_logic_vector(0 downto 0);
    signal cmp_2111 : std_logic_vector(0 downto 0);
    signal conv112_2157 : std_logic_vector(31 downto 0);
    signal conv115_1953 : std_logic_vector(31 downto 0);
    signal conv17_1894 : std_logic_vector(31 downto 0);
    signal conv65_2024 : std_logic_vector(63 downto 0);
    signal conv68_1941 : std_logic_vector(63 downto 0);
    signal conv70_2028 : std_logic_vector(63 downto 0);
    signal conv73_1945 : std_logic_vector(63 downto 0);
    signal conv75_2032 : std_logic_vector(63 downto 0);
    signal conv90_2100 : std_logic_vector(31 downto 0);
    signal conv94_1949 : std_logic_vector(31 downto 0);
    signal conv_1881 : std_logic_vector(31 downto 0);
    signal idxprom86_2085 : std_logic_vector(63 downto 0);
    signal idxprom_2062 : std_logic_vector(63 downto 0);
    signal inc110_2141 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2146 : std_logic_vector(15 downto 0);
    signal inc_2132 : std_logic_vector(15 downto 0);
    signal indvar_1962 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2195 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2183 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1983 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2177 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1976 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2153 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2170 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1969 : std_logic_vector(15 downto 0);
    signal mul54_2015 : std_logic_vector(15 downto 0);
    signal mul76_2037 : std_logic_vector(63 downto 0);
    signal mul78_2047 : std_logic_vector(63 downto 0);
    signal mul_2005 : std_logic_vector(15 downto 0);
    signal ptr_deref_2072_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2072_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2072_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2072_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2072_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2094_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2094_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2094_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2094_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2094_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2094_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1887 : std_logic_vector(31 downto 0);
    signal shr116132_1959 : std_logic_vector(31 downto 0);
    signal shr131_1915 : std_logic_vector(15 downto 0);
    signal shr81_2058 : std_logic_vector(31 downto 0);
    signal shr85_2079 : std_logic_vector(63 downto 0);
    signal sub48_2010 : std_logic_vector(15 downto 0);
    signal sub61_1937 : std_logic_vector(15 downto 0);
    signal sub62_2020 : std_logic_vector(15 downto 0);
    signal sub_1926 : std_logic_vector(15 downto 0);
    signal tmp1_1995 : std_logic_vector(31 downto 0);
    signal tmp83_2073 : std_logic_vector(63 downto 0);
    signal type_cast_1885_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1913_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1919_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1930_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1957_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1965_wire : std_logic_vector(31 downto 0);
    signal type_cast_1968_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1973_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1975_wire : std_logic_vector(15 downto 0);
    signal type_cast_1980_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1982_wire : std_logic_vector(15 downto 0);
    signal type_cast_1986_wire : std_logic_vector(15 downto 0);
    signal type_cast_1988_wire : std_logic_vector(15 downto 0);
    signal type_cast_1993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2056_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2077_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2083_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2104_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2122_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2130_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2150_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2173_wire : std_logic_vector(15 downto 0);
    signal type_cast_2176_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2180_wire : std_logic_vector(15 downto 0);
    signal type_cast_2182_wire : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire : std_logic_vector(15 downto 0);
    signal type_cast_2188_wire : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2201_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2067_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2067_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2067_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2067_resized_base_address <= "00000000000000";
    array_obj_ref_2090_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2090_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2090_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2090_resized_base_address <= "00000000000000";
    ptr_deref_2072_word_offset_0 <= "00000000000000";
    ptr_deref_2094_word_offset_0 <= "00000000000000";
    type_cast_1885_wire_constant <= "00000000000000000000000000010000";
    type_cast_1913_wire_constant <= "0000000000000010";
    type_cast_1919_wire_constant <= "1111111111111111";
    type_cast_1930_wire_constant <= "1111111111111111";
    type_cast_1957_wire_constant <= "00000000000000000000000000000001";
    type_cast_1968_wire_constant <= "00000000000000000000000000000000";
    type_cast_1973_wire_constant <= "0000000000000000";
    type_cast_1980_wire_constant <= "0000000000000000";
    type_cast_1993_wire_constant <= "00000000000000000000000000000100";
    type_cast_2056_wire_constant <= "00000000000000000000000000000010";
    type_cast_2077_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2083_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2104_wire_constant <= "00000000000000000000000000000100";
    type_cast_2122_wire_constant <= "0000000000000100";
    type_cast_2130_wire_constant <= "0000000000000001";
    type_cast_2150_wire_constant <= "0000000000000000";
    type_cast_2176_wire_constant <= "0000000000000000";
    type_cast_2193_wire_constant <= "00000000000000000000000000000001";
    type_cast_2201_wire_constant <= "0000000000000001";
    phi_stmt_1962: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1965_wire & type_cast_1968_wire_constant;
      req <= phi_stmt_1962_req_0 & phi_stmt_1962_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1962",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1962_ack_0,
          idata => idata,
          odata => indvar_1962,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1962
    phi_stmt_1969: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1973_wire_constant & type_cast_1975_wire;
      req <= phi_stmt_1969_req_0 & phi_stmt_1969_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1969",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1969_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1969,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1969
    phi_stmt_1976: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1980_wire_constant & type_cast_1982_wire;
      req <= phi_stmt_1976_req_0 & phi_stmt_1976_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1976",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1976_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1976,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1976
    phi_stmt_1983: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1986_wire & type_cast_1988_wire;
      req <= phi_stmt_1983_req_0 & phi_stmt_1983_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1983",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1983_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1983,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1983
    phi_stmt_2170: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2173_wire & type_cast_2176_wire_constant;
      req <= phi_stmt_2170_req_0 & phi_stmt_2170_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2170",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2170_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2170,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2170
    phi_stmt_2177: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2180_wire & type_cast_2182_wire;
      req <= phi_stmt_2177_req_0 & phi_stmt_2177_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2177",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2177_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2177,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2177
    phi_stmt_2183: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2186_wire & type_cast_2188_wire;
      req <= phi_stmt_2183_req_0 & phi_stmt_2183_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2183",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2183_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2183,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2183
    -- flow-through select operator MUX_2152_inst
    input_dim1x_x2_2153 <= type_cast_2150_wire_constant when (cmp106_2137(0) /=  '0') else inc_2132;
    addr_of_2068_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2068_final_reg_req_0;
      addr_of_2068_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2068_final_reg_req_1;
      addr_of_2068_final_reg_ack_1<= rack(0);
      addr_of_2068_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2068_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2067_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2091_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2091_final_reg_req_0;
      addr_of_2091_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2091_final_reg_req_1;
      addr_of_2091_final_reg_ack_1<= rack(0);
      addr_of_2091_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2091_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2090_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1880_inst_req_0;
      type_cast_1880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1880_inst_req_1;
      type_cast_1880_inst_ack_1<= rack(0);
      type_cast_1880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1893_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1893_inst_req_0;
      type_cast_1893_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1893_inst_req_1;
      type_cast_1893_inst_ack_1<= rack(0);
      type_cast_1893_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1893_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1890,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1940_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1940_inst_req_0;
      type_cast_1940_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1940_inst_req_1;
      type_cast_1940_inst_ack_1<= rack(0);
      type_cast_1940_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1940_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1941,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1944_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1944_inst_req_0;
      type_cast_1944_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1944_inst_req_1;
      type_cast_1944_inst_ack_1<= rack(0);
      type_cast_1944_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1944_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1945,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1948_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1948_inst_req_0;
      type_cast_1948_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1948_inst_req_1;
      type_cast_1948_inst_ack_1<= rack(0);
      type_cast_1948_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1948_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1949,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1952_inst_req_0;
      type_cast_1952_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1952_inst_req_1;
      type_cast_1952_inst_ack_1<= rack(0);
      type_cast_1952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1952_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1953,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1965_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1965_inst_req_0;
      type_cast_1965_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1965_inst_req_1;
      type_cast_1965_inst_ack_1<= rack(0);
      type_cast_1965_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1965_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2195,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1965_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1975_inst_req_0;
      type_cast_1975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1975_inst_req_1;
      type_cast_1975_inst_ack_1<= rack(0);
      type_cast_1975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1975_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1982_inst_req_0;
      type_cast_1982_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1982_inst_req_1;
      type_cast_1982_inst_ack_1<= rack(0);
      type_cast_1982_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1982_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1982_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1986_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1986_inst_req_0;
      type_cast_1986_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1986_inst_req_1;
      type_cast_1986_inst_ack_1<= rack(0);
      type_cast_1986_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1986_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1986_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1988_inst_req_0;
      type_cast_1988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1988_inst_req_1;
      type_cast_1988_inst_ack_1<= rack(0);
      type_cast_1988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1988_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1988_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2023_inst_req_0;
      type_cast_2023_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2023_inst_req_1;
      type_cast_2023_inst_ack_1<= rack(0);
      type_cast_2023_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2023_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1969,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2024,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2027_inst_req_0;
      type_cast_2027_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2027_inst_req_1;
      type_cast_2027_inst_ack_1<= rack(0);
      type_cast_2027_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2027_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2020,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2028,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2031_inst_req_0;
      type_cast_2031_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2031_inst_req_1;
      type_cast_2031_inst_ack_1<= rack(0);
      type_cast_2031_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2031_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2032,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2061_inst_req_0;
      type_cast_2061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2061_inst_req_1;
      type_cast_2061_inst_ack_1<= rack(0);
      type_cast_2061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2099_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2099_inst_req_0;
      type_cast_2099_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2099_inst_req_1;
      type_cast_2099_inst_ack_1<= rack(0);
      type_cast_2099_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2099_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1969,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2100,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2140_inst_req_0;
      type_cast_2140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2140_inst_req_1;
      type_cast_2140_inst_ack_1<= rack(0);
      type_cast_2140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2156_inst_req_0;
      type_cast_2156_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2156_inst_req_1;
      type_cast_2156_inst_ack_1<= rack(0);
      type_cast_2156_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2156_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2157,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2173_inst_req_0;
      type_cast_2173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2173_inst_req_1;
      type_cast_2173_inst_ack_1<= rack(0);
      type_cast_2173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2173_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1976,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2180_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2182_inst_req_0;
      type_cast_2182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2182_inst_req_1;
      type_cast_2182_inst_ack_1<= rack(0);
      type_cast_2182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2182_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2186_inst_req_0;
      type_cast_2186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2186_inst_req_1;
      type_cast_2186_inst_ack_1<= rack(0);
      type_cast_2186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2188_inst_req_0;
      type_cast_2188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2188_inst_req_1;
      type_cast_2188_inst_ack_1<= rack(0);
      type_cast_2188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2188_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2067_index_1_rename
    process(R_idxprom_2066_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2066_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2066_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2067_index_1_resize
    process(idxprom_2062) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2062;
      ov := iv(13 downto 0);
      R_idxprom_2066_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2067_root_address_inst
    process(array_obj_ref_2067_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2067_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2067_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2090_index_1_rename
    process(R_idxprom86_2089_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2089_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2089_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2090_index_1_resize
    process(idxprom86_2085) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2085;
      ov := iv(13 downto 0);
      R_idxprom86_2089_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2090_root_address_inst
    process(array_obj_ref_2090_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2090_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2090_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2072_addr_0
    process(ptr_deref_2072_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2072_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2072_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2072_base_resize
    process(arrayidx82_2069) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2069;
      ov := iv(13 downto 0);
      ptr_deref_2072_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2072_gather_scatter
    process(ptr_deref_2072_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2072_data_0;
      ov(63 downto 0) := iv;
      tmp83_2073 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2072_root_address_inst
    process(ptr_deref_2072_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2072_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2094_addr_0
    process(ptr_deref_2094_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2094_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2094_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2094_base_resize
    process(arrayidx87_2092) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2092;
      ov := iv(13 downto 0);
      ptr_deref_2094_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2094_gather_scatter
    process(tmp83_2073) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2073;
      ov(63 downto 0) := iv;
      ptr_deref_2094_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2094_root_address_inst
    process(ptr_deref_2094_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2094_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2094_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2112_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2111;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2112_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2112_branch_req_0,
          ack0 => if_stmt_2112_branch_ack_0,
          ack1 => if_stmt_2112_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2163_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2162;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2163_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2163_branch_req_0,
          ack0 => if_stmt_2163_branch_ack_0,
          ack1 => if_stmt_2163_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1920_inst
    process(call7_1862) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1862, type_cast_1919_wire_constant, tmp_var);
      add45_1921 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1931_inst
    process(call9_1865) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1865, type_cast_1930_wire_constant, tmp_var);
      add58_1932 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2009_inst
    process(sub_1926, mul_2005) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1926, mul_2005, tmp_var);
      sub48_2010 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2019_inst
    process(sub61_1937, mul54_2015) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1937, mul54_2015, tmp_var);
      sub62_2020 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2123_inst
    process(input_dim2x_x1_1969) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1969, type_cast_2122_wire_constant, tmp_var);
      add98_2124 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2131_inst
    process(input_dim1x_x1_1976) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1976, type_cast_2130_wire_constant, tmp_var);
      inc_2132 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2145_inst
    process(inc110_2141, input_dim0x_x2_1983) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2141, input_dim0x_x2_1983, tmp_var);
      inc110x_xinput_dim0x_x2_2146 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1999_inst
    process(add_1899, tmp1_1995) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1899, tmp1_1995, tmp_var);
      add_src_0x_x0_2000 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2105_inst
    process(conv90_2100) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2100, type_cast_2104_wire_constant, tmp_var);
      add91_2106 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2194_inst
    process(indvar_1962) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1962, type_cast_2193_wire_constant, tmp_var);
      indvarx_xnext_2195 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2041_inst
    process(mul76_2037, conv70_2028) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2037, conv70_2028, tmp_var);
      add77_2042 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2051_inst
    process(mul78_2047, conv65_2024) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2047, conv65_2024, tmp_var);
      add79_2052 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2084_inst
    process(shr85_2079) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2079, type_cast_2083_wire_constant, tmp_var);
      idxprom86_2085 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2136_inst
    process(inc_2132, call1_1853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2132, call1_1853, tmp_var);
      cmp106_2137 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2161_inst
    process(conv112_2157, shr116132_1959) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2157, shr116132_1959, tmp_var);
      cmp117_2162 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1914_inst
    process(call_1850) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1850, type_cast_1913_wire_constant, tmp_var);
      shr131_1915 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1958_inst
    process(conv115_1953) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1953, type_cast_1957_wire_constant, tmp_var);
      shr116132_1959 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2057_inst
    process(add_src_0x_x0_2000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2000, type_cast_2056_wire_constant, tmp_var);
      shr81_2058 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2078_inst
    process(add79_2052) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2052, type_cast_2077_wire_constant, tmp_var);
      shr85_2079 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2004_inst
    process(input_dim0x_x2_1983, call13_1871) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1983, call13_1871, tmp_var);
      mul_2005 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2014_inst
    process(input_dim1x_x1_1976, call13_1871) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1976, call13_1871, tmp_var);
      mul54_2015 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1994_inst
    process(indvar_1962) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1962, type_cast_1993_wire_constant, tmp_var);
      tmp1_1995 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2036_inst
    process(conv75_2032, conv73_1945) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2032, conv73_1945, tmp_var);
      mul76_2037 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2046_inst
    process(add77_2042, conv68_1941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2042, conv68_1941, tmp_var);
      mul78_2047 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1898_inst
    process(shl_1887, conv17_1894) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1887, conv17_1894, tmp_var);
      add_1899 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1886_inst
    process(conv_1881) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1881, type_cast_1885_wire_constant, tmp_var);
      shl_1887 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1925_inst
    process(add45_1921, call14_1874) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1921, call14_1874, tmp_var);
      sub_1926 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1936_inst
    process(add58_1932, call14_1874) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1932, call14_1874, tmp_var);
      sub61_1937 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2110_inst
    process(add91_2106, conv94_1949) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2106, conv94_1949, tmp_var);
      cmp_2111 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2067_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2066_scaled;
      array_obj_ref_2067_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2067_index_offset_req_0;
      array_obj_ref_2067_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2067_index_offset_req_1;
      array_obj_ref_2067_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2090_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2089_scaled;
      array_obj_ref_2090_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2090_index_offset_req_0;
      array_obj_ref_2090_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2090_index_offset_req_1;
      array_obj_ref_2090_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2072_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2072_load_0_req_0;
      ptr_deref_2072_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2072_load_0_req_1;
      ptr_deref_2072_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2072_word_address_0;
      ptr_deref_2072_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2094_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2094_store_0_req_0;
      ptr_deref_2094_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2094_store_0_req_1;
      ptr_deref_2094_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2094_word_address_0;
      data_in <= ptr_deref_2094_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1907_inst RPIPE_Block1_start_1904_inst RPIPE_Block1_start_1901_inst RPIPE_Block1_start_1889_inst RPIPE_Block1_start_1876_inst RPIPE_Block1_start_1873_inst RPIPE_Block1_start_1870_inst RPIPE_Block1_start_1867_inst RPIPE_Block1_start_1864_inst RPIPE_Block1_start_1861_inst RPIPE_Block1_start_1858_inst RPIPE_Block1_start_1855_inst RPIPE_Block1_start_1852_inst RPIPE_Block1_start_1849_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1907_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1904_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1901_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1889_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1876_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1873_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1870_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1867_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1864_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1861_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1858_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1855_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1852_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1849_inst_req_0;
      RPIPE_Block1_start_1907_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1904_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1901_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1889_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1876_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1873_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1870_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1867_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1864_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1861_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1858_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1855_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1852_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1849_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1907_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1904_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1901_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1889_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1876_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1873_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1870_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1867_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1864_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1861_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1858_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1855_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1852_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1849_inst_req_1;
      RPIPE_Block1_start_1907_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1904_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1901_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1889_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1876_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1873_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1870_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1867_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1864_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1861_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1858_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1855_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1852_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1849_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call22_1908 <= data_out(223 downto 208);
      call20_1905 <= data_out(207 downto 192);
      call18_1902 <= data_out(191 downto 176);
      call16_1890 <= data_out(175 downto 160);
      call15_1877 <= data_out(159 downto 144);
      call14_1874 <= data_out(143 downto 128);
      call13_1871 <= data_out(127 downto 112);
      call11_1868 <= data_out(111 downto 96);
      call9_1865 <= data_out(95 downto 80);
      call7_1862 <= data_out(79 downto 64);
      call5_1859 <= data_out(63 downto 48);
      call3_1856 <= data_out(47 downto 32);
      call1_1853 <= data_out(31 downto 16);
      call_1850 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2199_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2199_inst_req_0;
      WPIPE_Block1_done_2199_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2199_inst_req_1;
      WPIPE_Block1_done_2199_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2201_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5763_start: Boolean;
  signal convTransposeC_CP_5763_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2250_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2250_inst_ack_1 : boolean;
  signal type_cast_2305_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2228_inst_ack_1 : boolean;
  signal type_cast_2305_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2231_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2234_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2228_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2237_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2237_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2262_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2268_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2228_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2225_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2265_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2237_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2234_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2234_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2265_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2250_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2265_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2222_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2231_inst_ack_1 : boolean;
  signal type_cast_2254_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2225_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2234_inst_ack_1 : boolean;
  signal type_cast_2254_inst_ack_0 : boolean;
  signal type_cast_2241_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2262_inst_req_0 : boolean;
  signal type_cast_2254_inst_req_1 : boolean;
  signal type_cast_2254_inst_ack_1 : boolean;
  signal type_cast_2241_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2262_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2225_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2268_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2237_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2228_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_0 : boolean;
  signal type_cast_2301_inst_req_0 : boolean;
  signal type_cast_2305_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2225_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2262_inst_ack_1 : boolean;
  signal type_cast_2305_inst_req_0 : boolean;
  signal type_cast_2241_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2231_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2268_inst_ack_1 : boolean;
  signal type_cast_2241_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2231_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2250_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_ack_1 : boolean;
  signal type_cast_2301_inst_ack_0 : boolean;
  signal type_cast_2395_inst_ack_0 : boolean;
  signal type_cast_2395_inst_req_1 : boolean;
  signal type_cast_2309_inst_req_0 : boolean;
  signal type_cast_2313_inst_req_1 : boolean;
  signal type_cast_2313_inst_ack_1 : boolean;
  signal type_cast_2313_inst_ack_0 : boolean;
  signal type_cast_2313_inst_req_0 : boolean;
  signal type_cast_2395_inst_req_0 : boolean;
  signal type_cast_2301_inst_ack_1 : boolean;
  signal type_cast_2309_inst_req_1 : boolean;
  signal type_cast_2309_inst_ack_1 : boolean;
  signal type_cast_2301_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2268_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2265_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2210_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2210_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2210_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2210_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2213_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2213_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2213_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2213_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2219_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2219_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2219_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2219_inst_ack_1 : boolean;
  signal type_cast_2395_inst_ack_1 : boolean;
  signal type_cast_2399_inst_req_0 : boolean;
  signal type_cast_2399_inst_ack_0 : boolean;
  signal type_cast_2399_inst_req_1 : boolean;
  signal type_cast_2399_inst_ack_1 : boolean;
  signal type_cast_2403_inst_req_0 : boolean;
  signal type_cast_2403_inst_ack_0 : boolean;
  signal type_cast_2403_inst_req_1 : boolean;
  signal type_cast_2403_inst_ack_1 : boolean;
  signal type_cast_2433_inst_req_0 : boolean;
  signal type_cast_2433_inst_ack_0 : boolean;
  signal type_cast_2433_inst_req_1 : boolean;
  signal type_cast_2433_inst_ack_1 : boolean;
  signal array_obj_ref_2439_index_offset_req_0 : boolean;
  signal array_obj_ref_2439_index_offset_ack_0 : boolean;
  signal array_obj_ref_2439_index_offset_req_1 : boolean;
  signal array_obj_ref_2439_index_offset_ack_1 : boolean;
  signal addr_of_2440_final_reg_req_0 : boolean;
  signal addr_of_2440_final_reg_ack_0 : boolean;
  signal addr_of_2440_final_reg_req_1 : boolean;
  signal addr_of_2440_final_reg_ack_1 : boolean;
  signal ptr_deref_2444_load_0_req_0 : boolean;
  signal ptr_deref_2444_load_0_ack_0 : boolean;
  signal ptr_deref_2444_load_0_req_1 : boolean;
  signal ptr_deref_2444_load_0_ack_1 : boolean;
  signal array_obj_ref_2462_index_offset_req_0 : boolean;
  signal array_obj_ref_2462_index_offset_ack_0 : boolean;
  signal array_obj_ref_2462_index_offset_req_1 : boolean;
  signal array_obj_ref_2462_index_offset_ack_1 : boolean;
  signal addr_of_2463_final_reg_req_0 : boolean;
  signal addr_of_2463_final_reg_ack_0 : boolean;
  signal addr_of_2463_final_reg_req_1 : boolean;
  signal addr_of_2463_final_reg_ack_1 : boolean;
  signal ptr_deref_2466_store_0_req_0 : boolean;
  signal ptr_deref_2466_store_0_ack_0 : boolean;
  signal ptr_deref_2466_store_0_req_1 : boolean;
  signal ptr_deref_2466_store_0_ack_1 : boolean;
  signal type_cast_2471_inst_req_0 : boolean;
  signal type_cast_2471_inst_ack_0 : boolean;
  signal type_cast_2471_inst_req_1 : boolean;
  signal type_cast_2471_inst_ack_1 : boolean;
  signal if_stmt_2484_branch_req_0 : boolean;
  signal if_stmt_2484_branch_ack_1 : boolean;
  signal if_stmt_2484_branch_ack_0 : boolean;
  signal type_cast_2512_inst_req_0 : boolean;
  signal type_cast_2512_inst_ack_0 : boolean;
  signal type_cast_2512_inst_req_1 : boolean;
  signal type_cast_2512_inst_ack_1 : boolean;
  signal type_cast_2528_inst_req_0 : boolean;
  signal type_cast_2528_inst_ack_0 : boolean;
  signal type_cast_2528_inst_req_1 : boolean;
  signal type_cast_2528_inst_ack_1 : boolean;
  signal if_stmt_2535_branch_req_0 : boolean;
  signal if_stmt_2535_branch_ack_1 : boolean;
  signal if_stmt_2535_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2571_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2571_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2571_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2571_inst_ack_1 : boolean;
  signal phi_stmt_2334_req_0 : boolean;
  signal phi_stmt_2341_req_0 : boolean;
  signal phi_stmt_2348_req_1 : boolean;
  signal type_cast_2358_inst_req_0 : boolean;
  signal type_cast_2358_inst_ack_0 : boolean;
  signal type_cast_2358_inst_req_1 : boolean;
  signal type_cast_2358_inst_ack_1 : boolean;
  signal phi_stmt_2355_req_0 : boolean;
  signal type_cast_2340_inst_req_0 : boolean;
  signal type_cast_2340_inst_ack_0 : boolean;
  signal type_cast_2340_inst_req_1 : boolean;
  signal type_cast_2340_inst_ack_1 : boolean;
  signal phi_stmt_2334_req_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal phi_stmt_2341_req_1 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal phi_stmt_2348_req_0 : boolean;
  signal type_cast_2360_inst_req_0 : boolean;
  signal type_cast_2360_inst_ack_0 : boolean;
  signal type_cast_2360_inst_req_1 : boolean;
  signal type_cast_2360_inst_ack_1 : boolean;
  signal phi_stmt_2355_req_1 : boolean;
  signal phi_stmt_2334_ack_0 : boolean;
  signal phi_stmt_2341_ack_0 : boolean;
  signal phi_stmt_2348_ack_0 : boolean;
  signal phi_stmt_2355_ack_0 : boolean;
  signal phi_stmt_2542_req_1 : boolean;
  signal type_cast_2552_inst_req_0 : boolean;
  signal type_cast_2552_inst_ack_0 : boolean;
  signal type_cast_2552_inst_req_1 : boolean;
  signal type_cast_2552_inst_ack_1 : boolean;
  signal phi_stmt_2549_req_0 : boolean;
  signal type_cast_2558_inst_req_0 : boolean;
  signal type_cast_2558_inst_ack_0 : boolean;
  signal type_cast_2558_inst_req_1 : boolean;
  signal type_cast_2558_inst_ack_1 : boolean;
  signal phi_stmt_2555_req_0 : boolean;
  signal type_cast_2545_inst_req_0 : boolean;
  signal type_cast_2545_inst_ack_0 : boolean;
  signal type_cast_2545_inst_req_1 : boolean;
  signal type_cast_2545_inst_ack_1 : boolean;
  signal phi_stmt_2542_req_0 : boolean;
  signal type_cast_2554_inst_req_0 : boolean;
  signal type_cast_2554_inst_ack_0 : boolean;
  signal type_cast_2554_inst_req_1 : boolean;
  signal type_cast_2554_inst_ack_1 : boolean;
  signal phi_stmt_2549_req_1 : boolean;
  signal type_cast_2560_inst_req_0 : boolean;
  signal type_cast_2560_inst_ack_0 : boolean;
  signal type_cast_2560_inst_req_1 : boolean;
  signal type_cast_2560_inst_ack_1 : boolean;
  signal phi_stmt_2555_req_1 : boolean;
  signal phi_stmt_2542_ack_0 : boolean;
  signal phi_stmt_2549_ack_0 : boolean;
  signal phi_stmt_2555_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5763: Block -- control-path 
    signal convTransposeC_CP_5763_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5763_elements(0) <= convTransposeC_CP_5763_start;
    convTransposeC_CP_5763_symbol <= convTransposeC_CP_5763_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2208/$entry
      -- CP-element group 0: 	 branch_block_stmt_2208/branch_block_stmt_2208__entry__
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269__entry__
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/$entry
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Sample/rr
      -- 
    cr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => type_cast_2254_inst_req_1); -- 
    cr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => type_cast_2241_inst_req_1); -- 
    rr_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => RPIPE_Block2_start_2210_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2208/merge_stmt_2541__exit__
      -- CP-element group 1: 	 branch_block_stmt_2208/assign_stmt_2567__entry__
      -- CP-element group 1: 	 branch_block_stmt_2208/assign_stmt_2567__exit__
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2208/assign_stmt_2567/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/assign_stmt_2567/$exit
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Update/cr
      -- 
    rr_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2340_inst_req_0); -- 
    cr_6517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2340_inst_req_1); -- 
    rr_6535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2347_inst_req_0); -- 
    cr_6540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2347_inst_req_1); -- 
    rr_6558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2351_inst_req_0); -- 
    cr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2351_inst_req_1); -- 
    rr_6581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2360_inst_req_0); -- 
    cr_6586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2360_inst_req_1); -- 
    convTransposeC_CP_5763_elements(1) <= convTransposeC_CP_5763_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Update/cr
      -- 
    ra_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2210_inst_ack_0, ack => convTransposeC_CP_5763_elements(2)); -- 
    cr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(2), ack => RPIPE_Block2_start_2210_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2210_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Sample/rr
      -- 
    ca_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2210_inst_ack_1, ack => convTransposeC_CP_5763_elements(3)); -- 
    rr_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(3), ack => RPIPE_Block2_start_2213_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Update/cr
      -- 
    ra_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2213_inst_ack_0, ack => convTransposeC_CP_5763_elements(4)); -- 
    cr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(4), ack => RPIPE_Block2_start_2213_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2213_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Sample/rr
      -- 
    ca_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2213_inst_ack_1, ack => convTransposeC_CP_5763_elements(5)); -- 
    rr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(5), ack => RPIPE_Block2_start_2216_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Update/cr
      -- 
    ra_5840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_0, ack => convTransposeC_CP_5763_elements(6)); -- 
    cr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(6), ack => RPIPE_Block2_start_2216_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2216_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Sample/rr
      -- 
    ca_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_1, ack => convTransposeC_CP_5763_elements(7)); -- 
    rr_5853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(7), ack => RPIPE_Block2_start_2219_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Update/cr
      -- 
    ra_5854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2219_inst_ack_0, ack => convTransposeC_CP_5763_elements(8)); -- 
    cr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(8), ack => RPIPE_Block2_start_2219_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2219_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_sample_start_
      -- 
    ca_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2219_inst_ack_1, ack => convTransposeC_CP_5763_elements(9)); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(9), ack => RPIPE_Block2_start_2222_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_update_start_
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2222_inst_ack_0, ack => convTransposeC_CP_5763_elements(10)); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(10), ack => RPIPE_Block2_start_2222_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2222_update_completed_
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2222_inst_ack_1, ack => convTransposeC_CP_5763_elements(11)); -- 
    rr_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(11), ack => RPIPE_Block2_start_2225_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Sample/$exit
      -- 
    ra_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2225_inst_ack_0, ack => convTransposeC_CP_5763_elements(12)); -- 
    cr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(12), ack => RPIPE_Block2_start_2225_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2225_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Sample/$entry
      -- 
    ca_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2225_inst_ack_1, ack => convTransposeC_CP_5763_elements(13)); -- 
    rr_5895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(13), ack => RPIPE_Block2_start_2228_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_update_start_
      -- 
    ra_5896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2228_inst_ack_0, ack => convTransposeC_CP_5763_elements(14)); -- 
    cr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(14), ack => RPIPE_Block2_start_2228_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2228_update_completed_
      -- 
    ca_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2228_inst_ack_1, ack => convTransposeC_CP_5763_elements(15)); -- 
    rr_5909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(15), ack => RPIPE_Block2_start_2231_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Sample/ra
      -- 
    ra_5910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2231_inst_ack_0, ack => convTransposeC_CP_5763_elements(16)); -- 
    cr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(16), ack => RPIPE_Block2_start_2231_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2231_update_completed_
      -- 
    ca_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2231_inst_ack_1, ack => convTransposeC_CP_5763_elements(17)); -- 
    rr_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(17), ack => RPIPE_Block2_start_2234_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Sample/$exit
      -- 
    ra_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2234_inst_ack_0, ack => convTransposeC_CP_5763_elements(18)); -- 
    cr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(18), ack => RPIPE_Block2_start_2234_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2234_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Sample/$entry
      -- 
    ca_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2234_inst_ack_1, ack => convTransposeC_CP_5763_elements(19)); -- 
    rr_5937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(19), ack => RPIPE_Block2_start_2237_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Sample/$exit
      -- 
    ra_5938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2237_inst_ack_0, ack => convTransposeC_CP_5763_elements(20)); -- 
    cr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(20), ack => RPIPE_Block2_start_2237_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2237_update_completed_
      -- 
    ca_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2237_inst_ack_1, ack => convTransposeC_CP_5763_elements(21)); -- 
    rr_5951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(21), ack => type_cast_2241_inst_req_0); -- 
    rr_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(21), ack => RPIPE_Block2_start_2250_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Sample/ra
      -- 
    ra_5952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2241_inst_ack_0, ack => convTransposeC_CP_5763_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2241_Update/ca
      -- 
    ca_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2241_inst_ack_1, ack => convTransposeC_CP_5763_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Sample/ra
      -- 
    ra_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2250_inst_ack_0, ack => convTransposeC_CP_5763_elements(24)); -- 
    cr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(24), ack => RPIPE_Block2_start_2250_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2250_update_completed_
      -- 
    ca_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2250_inst_ack_1, ack => convTransposeC_CP_5763_elements(25)); -- 
    rr_5979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(25), ack => type_cast_2254_inst_req_0); -- 
    rr_5993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(25), ack => RPIPE_Block2_start_2262_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Sample/ra
      -- 
    ra_5980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_0, ack => convTransposeC_CP_5763_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/type_cast_2254_Update/ca
      -- 
    ca_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_1, ack => convTransposeC_CP_5763_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_update_start_
      -- 
    ra_5994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2262_inst_ack_0, ack => convTransposeC_CP_5763_elements(28)); -- 
    cr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(28), ack => RPIPE_Block2_start_2262_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2262_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_sample_start_
      -- 
    ca_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2262_inst_ack_1, ack => convTransposeC_CP_5763_elements(29)); -- 
    rr_6007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(29), ack => RPIPE_Block2_start_2265_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Sample/ra
      -- 
    ra_6008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2265_inst_ack_0, ack => convTransposeC_CP_5763_elements(30)); -- 
    cr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(30), ack => RPIPE_Block2_start_2265_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2265_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Sample/rr
      -- 
    ca_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2265_inst_ack_1, ack => convTransposeC_CP_5763_elements(31)); -- 
    rr_6021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(31), ack => RPIPE_Block2_start_2268_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Sample/$exit
      -- 
    ra_6022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2268_inst_ack_0, ack => convTransposeC_CP_5763_elements(32)); -- 
    cr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(32), ack => RPIPE_Block2_start_2268_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/RPIPE_Block2_start_2268_Update/ca
      -- 
    ca_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2268_inst_ack_1, ack => convTransposeC_CP_5763_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269__exit__
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331__entry__
      -- CP-element group 34: 	 branch_block_stmt_2208/assign_stmt_2211_to_assign_stmt_2269/$exit
      -- 
    cr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2305_inst_req_1); -- 
    rr_6038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2301_inst_req_0); -- 
    rr_6052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2305_inst_req_0); -- 
    rr_6066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2309_inst_req_0); -- 
    cr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2313_inst_req_1); -- 
    rr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2313_inst_req_0); -- 
    cr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2309_inst_req_1); -- 
    cr_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2301_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(23) & convTransposeC_CP_5763_elements(27) & convTransposeC_CP_5763_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Sample/ra
      -- 
    ra_6039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2301_inst_ack_0, ack => convTransposeC_CP_5763_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2301_Update/$exit
      -- 
    ca_6044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2301_inst_ack_1, ack => convTransposeC_CP_5763_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_sample_completed_
      -- 
    ra_6053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_0, ack => convTransposeC_CP_5763_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2305_update_completed_
      -- 
    ca_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_1, ack => convTransposeC_CP_5763_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_sample_completed_
      -- 
    ra_6067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_0, ack => convTransposeC_CP_5763_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2309_Update/ca
      -- 
    ca_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2309_inst_ack_1, ack => convTransposeC_CP_5763_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_sample_completed_
      -- 
    ra_6081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2313_inst_ack_0, ack => convTransposeC_CP_5763_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/type_cast_2313_update_completed_
      -- 
    ca_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2313_inst_ack_1, ack => convTransposeC_CP_5763_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331/$exit
      -- CP-element group 43: 	 branch_block_stmt_2208/assign_stmt_2276_to_assign_stmt_2331__exit__
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/cr
      -- 
    rr_6486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(43), ack => type_cast_2358_inst_req_0); -- 
    cr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(43), ack => type_cast_2358_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(36) & convTransposeC_CP_5763_elements(38) & convTransposeC_CP_5763_elements(40) & convTransposeC_CP_5763_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Sample/$exit
      -- 
    ra_6098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_0, ack => convTransposeC_CP_5763_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Update/ca
      -- 
    ca_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2395_inst_ack_1, ack => convTransposeC_CP_5763_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Sample/ra
      -- 
    ra_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_0, ack => convTransposeC_CP_5763_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Update/ca
      -- 
    ca_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_1, ack => convTransposeC_CP_5763_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Sample/ra
      -- 
    ra_6126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_0, ack => convTransposeC_CP_5763_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Update/ca
      -- 
    ca_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_1, ack => convTransposeC_CP_5763_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Sample/ra
      -- 
    ra_6140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_0, ack => convTransposeC_CP_5763_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Sample/req
      -- 
    ca_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_1, ack => convTransposeC_CP_5763_elements(51)); -- 
    req_6170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(51), ack => array_obj_ref_2439_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Sample/ack
      -- 
    ack_6171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2439_index_offset_ack_0, ack => convTransposeC_CP_5763_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_request/req
      -- 
    ack_6176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2439_index_offset_ack_1, ack => convTransposeC_CP_5763_elements(53)); -- 
    req_6185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(53), ack => addr_of_2440_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_request/ack
      -- 
    ack_6186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2440_final_reg_ack_0, ack => convTransposeC_CP_5763_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/word_0/rr
      -- 
    ack_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2440_final_reg_ack_1, ack => convTransposeC_CP_5763_elements(55)); -- 
    rr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(55), ack => ptr_deref_2444_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Sample/word_access_start/word_0/ra
      -- 
    ra_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2444_load_0_ack_0, ack => convTransposeC_CP_5763_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/ptr_deref_2444_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/ptr_deref_2444_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/ptr_deref_2444_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/ptr_deref_2444_Merge/merge_ack
      -- 
    ca_6236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2444_load_0_ack_1, ack => convTransposeC_CP_5763_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Sample/req
      -- 
    req_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(58), ack => array_obj_ref_2462_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(45) & convTransposeC_CP_5763_elements(47) & convTransposeC_CP_5763_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Sample/ack
      -- 
    ack_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2462_index_offset_ack_0, ack => convTransposeC_CP_5763_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_request/req
      -- 
    ack_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2462_index_offset_ack_1, ack => convTransposeC_CP_5763_elements(60)); -- 
    req_6281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(60), ack => addr_of_2463_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_request/ack
      -- 
    ack_6282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2463_final_reg_ack_0, ack => convTransposeC_CP_5763_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_word_addrgen/root_register_ack
      -- 
    ack_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2463_final_reg_ack_1, ack => convTransposeC_CP_5763_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/ptr_deref_2466_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/ptr_deref_2466_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/ptr_deref_2466_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/ptr_deref_2466_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/word_0/rr
      -- 
    rr_6325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(63), ack => ptr_deref_2466_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(57) & convTransposeC_CP_5763_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Sample/word_access_start/word_0/ra
      -- 
    ra_6326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2466_store_0_ack_0, ack => convTransposeC_CP_5763_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/word_0/ca
      -- 
    ca_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2466_store_0_ack_1, ack => convTransposeC_CP_5763_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Sample/ra
      -- 
    ra_6346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_0, ack => convTransposeC_CP_5763_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Update/ca
      -- 
    ca_6351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2471_inst_ack_1, ack => convTransposeC_CP_5763_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/$exit
      -- CP-element group 68: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483__exit__
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484__entry__
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2208/R_cmp_2485_place
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2208/if_stmt_2484_else_link/$entry
      -- 
    branch_req_6359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(68), ack => if_stmt_2484_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(52) & convTransposeC_CP_5763_elements(59) & convTransposeC_CP_5763_elements(65) & convTransposeC_CP_5763_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2208/merge_stmt_2490__exit__
      -- CP-element group 69: 	 branch_block_stmt_2208/assign_stmt_2496__entry__
      -- CP-element group 69: 	 branch_block_stmt_2208/assign_stmt_2496__exit__
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2208/if_stmt_2484_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2208/if_stmt_2484_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2208/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2208/assign_stmt_2496/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/assign_stmt_2496/$exit
      -- CP-element group 69: 	 branch_block_stmt_2208/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2208/merge_stmt_2490_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2208/merge_stmt_2490_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/merge_stmt_2490_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2208/merge_stmt_2490_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2484_branch_ack_1, ack => convTransposeC_CP_5763_elements(69)); -- 
    rr_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2545_inst_req_0); -- 
    cr_6701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2545_inst_req_1); -- 
    rr_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2554_inst_req_0); -- 
    cr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2554_inst_req_1); -- 
    rr_6742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2560_inst_req_0); -- 
    cr_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2560_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2208/merge_stmt_2498__exit__
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534__entry__
      -- CP-element group 70: 	 branch_block_stmt_2208/if_stmt_2484_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2208/if_stmt_2484_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2208/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2208/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2208/merge_stmt_2498_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2208/merge_stmt_2498_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2208/merge_stmt_2498_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2208/merge_stmt_2498_PhiAck/dummy
      -- 
    else_choice_transition_6368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2484_branch_ack_0, ack => convTransposeC_CP_5763_elements(70)); -- 
    rr_6384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2512_inst_req_0); -- 
    cr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2512_inst_req_1); -- 
    cr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2528_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Sample/ra
      -- 
    ra_6385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_0, ack => convTransposeC_CP_5763_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2512_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Sample/rr
      -- 
    ca_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_1, ack => convTransposeC_CP_5763_elements(72)); -- 
    rr_6398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(72), ack => type_cast_2528_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Sample/ra
      -- 
    ra_6399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2528_inst_ack_0, ack => convTransposeC_CP_5763_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534__exit__
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535__entry__
      -- CP-element group 74: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/$exit
      -- CP-element group 74: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2208/assign_stmt_2504_to_assign_stmt_2534/type_cast_2528_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2208/R_cmp122_2536_place
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2208/if_stmt_2535_else_link/$entry
      -- 
    ca_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2528_inst_ack_1, ack => convTransposeC_CP_5763_elements(74)); -- 
    branch_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(74), ack => if_stmt_2535_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2208/merge_stmt_2569__exit__
      -- CP-element group 75: 	 branch_block_stmt_2208/assign_stmt_2574__entry__
      -- CP-element group 75: 	 branch_block_stmt_2208/if_stmt_2535_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2208/if_stmt_2535_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2208/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2208/assign_stmt_2574/$entry
      -- CP-element group 75: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2208/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2208/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2208/merge_stmt_2569_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2208/merge_stmt_2569_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2208/merge_stmt_2569_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2208/merge_stmt_2569_PhiAck/dummy
      -- 
    if_choice_transition_6417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2535_branch_ack_1, ack => convTransposeC_CP_5763_elements(75)); -- 
    req_6437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(75), ack => WPIPE_Block2_done_2571_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2208/if_stmt_2535_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2208/if_stmt_2535_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2535_branch_ack_0, ack => convTransposeC_CP_5763_elements(76)); -- 
    rr_6647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2552_inst_req_0); -- 
    cr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2552_inst_req_1); -- 
    rr_6670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2558_inst_req_0); -- 
    cr_6675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2558_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Update/req
      -- 
    ack_6438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2571_inst_ack_0, ack => convTransposeC_CP_5763_elements(77)); -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(77), ack => WPIPE_Block2_done_2571_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2208/$exit
      -- CP-element group 78: 	 branch_block_stmt_2208/branch_block_stmt_2208__exit__
      -- CP-element group 78: 	 branch_block_stmt_2208/assign_stmt_2574__exit__
      -- CP-element group 78: 	 branch_block_stmt_2208/return__
      -- CP-element group 78: 	 branch_block_stmt_2208/merge_stmt_2576__exit__
      -- CP-element group 78: 	 branch_block_stmt_2208/assign_stmt_2574/$exit
      -- CP-element group 78: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2208/assign_stmt_2574/WPIPE_Block2_done_2571_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2208/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2208/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2208/merge_stmt_2576_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2208/merge_stmt_2576_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2208/merge_stmt_2576_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2208/merge_stmt_2576_PhiAck/dummy
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2571_inst_ack_1, ack => convTransposeC_CP_5763_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/$exit
      -- CP-element group 79: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2338_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_req
      -- 
    phi_stmt_2334_req_6454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2334_req_6454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(79), ack => phi_stmt_2334_req_0); -- 
    -- Element group convTransposeC_CP_5763_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/$exit
      -- CP-element group 80: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2345_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_req
      -- 
    phi_stmt_2341_req_6462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2341_req_6462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(80), ack => phi_stmt_2341_req_0); -- 
    -- Element group convTransposeC_CP_5763_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/$exit
      -- CP-element group 81: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2354_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_req
      -- 
    phi_stmt_2348_req_6470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2348_req_6470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(81), ack => phi_stmt_2348_req_1); -- 
    -- Element group convTransposeC_CP_5763_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Sample/ra
      -- 
    ra_6487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_0, ack => convTransposeC_CP_5763_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/Update/ca
      -- 
    ca_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_1, ack => convTransposeC_CP_5763_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/$exit
      -- CP-element group 84: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/$exit
      -- CP-element group 84: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2358/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_req
      -- 
    phi_stmt_2355_req_6493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2355_req_6493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(84), ack => phi_stmt_2355_req_0); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(82) & convTransposeC_CP_5763_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2208/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(79) & convTransposeC_CP_5763_elements(80) & convTransposeC_CP_5763_elements(81) & convTransposeC_CP_5763_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Sample/ra
      -- 
    ra_6513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2340_inst_ack_0, ack => convTransposeC_CP_5763_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/Update/ca
      -- 
    ca_6518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2340_inst_ack_1, ack => convTransposeC_CP_5763_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/$exit
      -- CP-element group 88: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/$exit
      -- CP-element group 88: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_sources/type_cast_2340/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2334/phi_stmt_2334_req
      -- 
    phi_stmt_2334_req_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2334_req_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(88), ack => phi_stmt_2334_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(86) & convTransposeC_CP_5763_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Sample/ra
      -- 
    ra_6536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => convTransposeC_CP_5763_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/Update/ca
      -- 
    ca_6541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => convTransposeC_CP_5763_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/$exit
      -- CP-element group 91: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/$exit
      -- CP-element group 91: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_sources/type_cast_2347/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2341/phi_stmt_2341_req
      -- 
    phi_stmt_2341_req_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2341_req_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(91), ack => phi_stmt_2341_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(89) & convTransposeC_CP_5763_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Sample/ra
      -- 
    ra_6559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convTransposeC_CP_5763_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/Update/ca
      -- 
    ca_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convTransposeC_CP_5763_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/$exit
      -- CP-element group 94: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/$exit
      -- CP-element group 94: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_sources/type_cast_2351/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2348/phi_stmt_2348_req
      -- 
    phi_stmt_2348_req_6565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2348_req_6565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(94), ack => phi_stmt_2348_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(92) & convTransposeC_CP_5763_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Sample/ra
      -- 
    ra_6582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2360_inst_ack_0, ack => convTransposeC_CP_5763_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/Update/ca
      -- 
    ca_6587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2360_inst_ack_1, ack => convTransposeC_CP_5763_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/$exit
      -- CP-element group 97: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/$exit
      -- CP-element group 97: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_sources/type_cast_2360/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2355/phi_stmt_2355_req
      -- 
    phi_stmt_2355_req_6588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2355_req_6588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(97), ack => phi_stmt_2355_req_1); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(95) & convTransposeC_CP_5763_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2208/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(88) & convTransposeC_CP_5763_elements(91) & convTransposeC_CP_5763_elements(94) & convTransposeC_CP_5763_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2208/merge_stmt_2333_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/$entry
      -- 
    convTransposeC_CP_5763_elements(99) <= OrReduce(convTransposeC_CP_5763_elements(85) & convTransposeC_CP_5763_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/phi_stmt_2334_ack
      -- 
    phi_stmt_2334_ack_6593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2334_ack_0, ack => convTransposeC_CP_5763_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/phi_stmt_2341_ack
      -- 
    phi_stmt_2341_ack_6594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2341_ack_0, ack => convTransposeC_CP_5763_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/phi_stmt_2348_ack
      -- 
    phi_stmt_2348_ack_6595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2348_ack_0, ack => convTransposeC_CP_5763_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/phi_stmt_2355_ack
      -- 
    phi_stmt_2355_ack_6596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2355_ack_0, ack => convTransposeC_CP_5763_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2395_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2208/merge_stmt_2333__exit__
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483__entry__
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2399_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2403_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2433_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2439_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2440_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2444_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/array_obj_ref_2462_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/addr_of_2463_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/ptr_deref_2466_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2208/assign_stmt_2367_to_assign_stmt_2483/type_cast_2471_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2208/merge_stmt_2333_PhiAck/$exit
      -- 
    cr_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2395_inst_req_1); -- 
    rr_6097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2395_inst_req_0); -- 
    rr_6111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2399_inst_req_0); -- 
    cr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2399_inst_req_1); -- 
    rr_6125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2403_inst_req_0); -- 
    cr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2403_inst_req_1); -- 
    rr_6139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2433_inst_req_0); -- 
    cr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2433_inst_req_1); -- 
    req_6175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => array_obj_ref_2439_index_offset_req_1); -- 
    req_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => addr_of_2440_final_reg_req_1); -- 
    cr_6235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => ptr_deref_2444_load_0_req_1); -- 
    req_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => array_obj_ref_2462_index_offset_req_1); -- 
    req_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => addr_of_2463_final_reg_req_1); -- 
    cr_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => ptr_deref_2466_store_0_req_1); -- 
    rr_6345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2471_inst_req_0); -- 
    cr_6350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2471_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(100) & convTransposeC_CP_5763_elements(101) & convTransposeC_CP_5763_elements(102) & convTransposeC_CP_5763_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/$exit
      -- CP-element group 105: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2548_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_req
      -- 
    phi_stmt_2542_req_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2542_req_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(105), ack => phi_stmt_2542_req_1); -- 
    -- Element group convTransposeC_CP_5763_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(76), ack => convTransposeC_CP_5763_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Sample/ra
      -- 
    ra_6648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2552_inst_ack_0, ack => convTransposeC_CP_5763_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/Update/ca
      -- 
    ca_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2552_inst_ack_1, ack => convTransposeC_CP_5763_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/$exit
      -- CP-element group 108: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/$exit
      -- CP-element group 108: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2552/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_req
      -- 
    phi_stmt_2549_req_6654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2549_req_6654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(108), ack => phi_stmt_2549_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(106) & convTransposeC_CP_5763_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/ra
      -- 
    ra_6671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2558_inst_ack_0, ack => convTransposeC_CP_5763_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/ca
      -- 
    ca_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2558_inst_ack_1, ack => convTransposeC_CP_5763_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/$exit
      -- CP-element group 111: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/$exit
      -- CP-element group 111: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_req
      -- 
    phi_stmt_2555_req_6677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2555_req_6677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(111), ack => phi_stmt_2555_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(109) & convTransposeC_CP_5763_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2208/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(105) & convTransposeC_CP_5763_elements(108) & convTransposeC_CP_5763_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Sample/ra
      -- 
    ra_6697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_0, ack => convTransposeC_CP_5763_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/Update/ca
      -- 
    ca_6702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_1, ack => convTransposeC_CP_5763_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/$exit
      -- CP-element group 115: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/$exit
      -- CP-element group 115: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_sources/type_cast_2545/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2542/phi_stmt_2542_req
      -- 
    phi_stmt_2542_req_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2542_req_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(115), ack => phi_stmt_2542_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(113) & convTransposeC_CP_5763_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Sample/ra
      -- 
    ra_6720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2554_inst_ack_0, ack => convTransposeC_CP_5763_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/Update/ca
      -- 
    ca_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2554_inst_ack_1, ack => convTransposeC_CP_5763_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/$exit
      -- CP-element group 118: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/$exit
      -- CP-element group 118: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_sources/type_cast_2554/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2549/phi_stmt_2549_req
      -- 
    phi_stmt_2549_req_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2549_req_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(118), ack => phi_stmt_2549_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(116) & convTransposeC_CP_5763_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/ra
      -- 
    ra_6743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_0, ack => convTransposeC_CP_5763_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/ca
      -- 
    ca_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_1, ack => convTransposeC_CP_5763_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/$exit
      -- CP-element group 121: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/$exit
      -- CP-element group 121: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_req
      -- 
    phi_stmt_2555_req_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2555_req_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(121), ack => phi_stmt_2555_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(119) & convTransposeC_CP_5763_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2208/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(115) & convTransposeC_CP_5763_elements(118) & convTransposeC_CP_5763_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2208/merge_stmt_2541_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2208/merge_stmt_2541_PhiAck/$entry
      -- 
    convTransposeC_CP_5763_elements(123) <= OrReduce(convTransposeC_CP_5763_elements(112) & convTransposeC_CP_5763_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2208/merge_stmt_2541_PhiAck/phi_stmt_2542_ack
      -- 
    phi_stmt_2542_ack_6754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2542_ack_0, ack => convTransposeC_CP_5763_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2208/merge_stmt_2541_PhiAck/phi_stmt_2549_ack
      -- 
    phi_stmt_2549_ack_6755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2549_ack_0, ack => convTransposeC_CP_5763_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2208/merge_stmt_2541_PhiAck/phi_stmt_2555_ack
      -- 
    phi_stmt_2555_ack_6756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2555_ack_0, ack => convTransposeC_CP_5763_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2208/merge_stmt_2541_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(124) & convTransposeC_CP_5763_elements(125) & convTransposeC_CP_5763_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2461_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2461_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2438_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2438_scaled : std_logic_vector(13 downto 0);
    signal add121_2331 : std_logic_vector(31 downto 0);
    signal add45_2282 : std_logic_vector(15 downto 0);
    signal add58_2293 : std_logic_vector(15 downto 0);
    signal add77_2414 : std_logic_vector(63 downto 0);
    signal add79_2424 : std_logic_vector(63 downto 0);
    signal add91_2478 : std_logic_vector(31 downto 0);
    signal add98_2496 : std_logic_vector(15 downto 0);
    signal add_2260 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2372 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2439_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2439_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2439_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2439_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2439_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2439_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2462_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2441 : std_logic_vector(31 downto 0);
    signal arrayidx87_2464 : std_logic_vector(31 downto 0);
    signal call11_2229 : std_logic_vector(15 downto 0);
    signal call13_2232 : std_logic_vector(15 downto 0);
    signal call14_2235 : std_logic_vector(15 downto 0);
    signal call15_2238 : std_logic_vector(15 downto 0);
    signal call16_2251 : std_logic_vector(15 downto 0);
    signal call18_2263 : std_logic_vector(15 downto 0);
    signal call1_2214 : std_logic_vector(15 downto 0);
    signal call20_2266 : std_logic_vector(15 downto 0);
    signal call22_2269 : std_logic_vector(15 downto 0);
    signal call3_2217 : std_logic_vector(15 downto 0);
    signal call5_2220 : std_logic_vector(15 downto 0);
    signal call7_2223 : std_logic_vector(15 downto 0);
    signal call9_2226 : std_logic_vector(15 downto 0);
    signal call_2211 : std_logic_vector(15 downto 0);
    signal cmp106_2509 : std_logic_vector(0 downto 0);
    signal cmp122_2534 : std_logic_vector(0 downto 0);
    signal cmp_2483 : std_logic_vector(0 downto 0);
    signal conv112_2529 : std_logic_vector(31 downto 0);
    signal conv115_2314 : std_logic_vector(31 downto 0);
    signal conv17_2255 : std_logic_vector(31 downto 0);
    signal conv65_2396 : std_logic_vector(63 downto 0);
    signal conv68_2302 : std_logic_vector(63 downto 0);
    signal conv70_2400 : std_logic_vector(63 downto 0);
    signal conv73_2306 : std_logic_vector(63 downto 0);
    signal conv75_2404 : std_logic_vector(63 downto 0);
    signal conv90_2472 : std_logic_vector(31 downto 0);
    signal conv94_2310 : std_logic_vector(31 downto 0);
    signal conv_2242 : std_logic_vector(31 downto 0);
    signal idxprom86_2457 : std_logic_vector(63 downto 0);
    signal idxprom_2434 : std_logic_vector(63 downto 0);
    signal inc110_2513 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2518 : std_logic_vector(15 downto 0);
    signal inc_2504 : std_logic_vector(15 downto 0);
    signal indvar_2334 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2567 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2555 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2355 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2549 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2348 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2525 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2542 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2341 : std_logic_vector(15 downto 0);
    signal mul54_2387 : std_logic_vector(15 downto 0);
    signal mul76_2409 : std_logic_vector(63 downto 0);
    signal mul78_2419 : std_logic_vector(63 downto 0);
    signal mul_2377 : std_logic_vector(15 downto 0);
    signal ptr_deref_2444_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2444_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2444_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2444_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2444_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2466_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2466_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2466_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2466_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2466_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2466_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2248 : std_logic_vector(31 downto 0);
    signal shr116137_2320 : std_logic_vector(31 downto 0);
    signal shr120138_2326 : std_logic_vector(31 downto 0);
    signal shr136_2276 : std_logic_vector(15 downto 0);
    signal shr81_2430 : std_logic_vector(31 downto 0);
    signal shr85_2451 : std_logic_vector(63 downto 0);
    signal sub48_2382 : std_logic_vector(15 downto 0);
    signal sub61_2298 : std_logic_vector(15 downto 0);
    signal sub62_2392 : std_logic_vector(15 downto 0);
    signal sub_2287 : std_logic_vector(15 downto 0);
    signal tmp1_2367 : std_logic_vector(31 downto 0);
    signal tmp83_2445 : std_logic_vector(63 downto 0);
    signal type_cast_2246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2274_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2280_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2291_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2318_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2324_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2338_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2340_wire : std_logic_vector(31 downto 0);
    signal type_cast_2345_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2347_wire : std_logic_vector(15 downto 0);
    signal type_cast_2351_wire : std_logic_vector(15 downto 0);
    signal type_cast_2354_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2358_wire : std_logic_vector(15 downto 0);
    signal type_cast_2360_wire : std_logic_vector(15 downto 0);
    signal type_cast_2365_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2449_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2476_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2494_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2502_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2522_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2545_wire : std_logic_vector(15 downto 0);
    signal type_cast_2548_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2552_wire : std_logic_vector(15 downto 0);
    signal type_cast_2554_wire : std_logic_vector(15 downto 0);
    signal type_cast_2558_wire : std_logic_vector(15 downto 0);
    signal type_cast_2560_wire : std_logic_vector(15 downto 0);
    signal type_cast_2565_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2573_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2439_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2439_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2439_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2439_resized_base_address <= "00000000000000";
    array_obj_ref_2462_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2462_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2462_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2462_resized_base_address <= "00000000000000";
    ptr_deref_2444_word_offset_0 <= "00000000000000";
    ptr_deref_2466_word_offset_0 <= "00000000000000";
    type_cast_2246_wire_constant <= "00000000000000000000000000010000";
    type_cast_2274_wire_constant <= "0000000000000001";
    type_cast_2280_wire_constant <= "1111111111111111";
    type_cast_2291_wire_constant <= "1111111111111111";
    type_cast_2318_wire_constant <= "00000000000000000000000000000010";
    type_cast_2324_wire_constant <= "00000000000000000000000000000001";
    type_cast_2338_wire_constant <= "00000000000000000000000000000000";
    type_cast_2345_wire_constant <= "0000000000000000";
    type_cast_2354_wire_constant <= "0000000000000000";
    type_cast_2365_wire_constant <= "00000000000000000000000000000100";
    type_cast_2428_wire_constant <= "00000000000000000000000000000010";
    type_cast_2449_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2455_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2476_wire_constant <= "00000000000000000000000000000100";
    type_cast_2494_wire_constant <= "0000000000000100";
    type_cast_2502_wire_constant <= "0000000000000001";
    type_cast_2522_wire_constant <= "0000000000000000";
    type_cast_2548_wire_constant <= "0000000000000000";
    type_cast_2565_wire_constant <= "00000000000000000000000000000001";
    type_cast_2573_wire_constant <= "0000000000000001";
    phi_stmt_2334: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2338_wire_constant & type_cast_2340_wire;
      req <= phi_stmt_2334_req_0 & phi_stmt_2334_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2334",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2334_ack_0,
          idata => idata,
          odata => indvar_2334,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2334
    phi_stmt_2341: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2345_wire_constant & type_cast_2347_wire;
      req <= phi_stmt_2341_req_0 & phi_stmt_2341_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2341",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2341_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2341,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2341
    phi_stmt_2348: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2351_wire & type_cast_2354_wire_constant;
      req <= phi_stmt_2348_req_0 & phi_stmt_2348_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2348",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2348_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2348,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2348
    phi_stmt_2355: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2358_wire & type_cast_2360_wire;
      req <= phi_stmt_2355_req_0 & phi_stmt_2355_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2355",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2355_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2355,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2355
    phi_stmt_2542: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2545_wire & type_cast_2548_wire_constant;
      req <= phi_stmt_2542_req_0 & phi_stmt_2542_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2542",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2542_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2542,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2542
    phi_stmt_2549: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2552_wire & type_cast_2554_wire;
      req <= phi_stmt_2549_req_0 & phi_stmt_2549_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2549",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2549_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2549,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2549
    phi_stmt_2555: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2558_wire & type_cast_2560_wire;
      req <= phi_stmt_2555_req_0 & phi_stmt_2555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2555",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2555_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2555
    -- flow-through select operator MUX_2524_inst
    input_dim1x_x2_2525 <= type_cast_2522_wire_constant when (cmp106_2509(0) /=  '0') else inc_2504;
    addr_of_2440_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2440_final_reg_req_0;
      addr_of_2440_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2440_final_reg_req_1;
      addr_of_2440_final_reg_ack_1<= rack(0);
      addr_of_2440_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2440_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2439_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2441,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2463_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2463_final_reg_req_0;
      addr_of_2463_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2463_final_reg_req_1;
      addr_of_2463_final_reg_ack_1<= rack(0);
      addr_of_2463_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2463_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2462_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2241_inst_req_0;
      type_cast_2241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2241_inst_req_1;
      type_cast_2241_inst_ack_1<= rack(0);
      type_cast_2241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2254_inst_req_0;
      type_cast_2254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2254_inst_req_1;
      type_cast_2254_inst_ack_1<= rack(0);
      type_cast_2254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2301_inst_req_0;
      type_cast_2301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2301_inst_req_1;
      type_cast_2301_inst_ack_1<= rack(0);
      type_cast_2301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2305_inst_req_0;
      type_cast_2305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2305_inst_req_1;
      type_cast_2305_inst_ack_1<= rack(0);
      type_cast_2305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2266,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2309_inst_req_0;
      type_cast_2309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2309_inst_req_1;
      type_cast_2309_inst_ack_1<= rack(0);
      type_cast_2309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2313_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2313_inst_req_0;
      type_cast_2313_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2313_inst_req_1;
      type_cast_2313_inst_ack_1<= rack(0);
      type_cast_2313_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2313_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2314,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2340_inst_req_0;
      type_cast_2340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2340_inst_req_1;
      type_cast_2340_inst_ack_1<= rack(0);
      type_cast_2340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2340_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2542,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2347_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2549,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2351_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2358_inst_req_0;
      type_cast_2358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2358_inst_req_1;
      type_cast_2358_inst_ack_1<= rack(0);
      type_cast_2358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2358_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2360_inst_req_0;
      type_cast_2360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2360_inst_req_1;
      type_cast_2360_inst_ack_1<= rack(0);
      type_cast_2360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2360_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2395_inst_req_0;
      type_cast_2395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2395_inst_req_1;
      type_cast_2395_inst_ack_1<= rack(0);
      type_cast_2395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2399_inst_req_0;
      type_cast_2399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2399_inst_req_1;
      type_cast_2399_inst_ack_1<= rack(0);
      type_cast_2399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2403_inst_req_0;
      type_cast_2403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2403_inst_req_1;
      type_cast_2403_inst_ack_1<= rack(0);
      type_cast_2403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2433_inst_req_0;
      type_cast_2433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2433_inst_req_1;
      type_cast_2433_inst_ack_1<= rack(0);
      type_cast_2433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2434,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2471_inst_req_0;
      type_cast_2471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2471_inst_req_1;
      type_cast_2471_inst_ack_1<= rack(0);
      type_cast_2471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2512_inst_req_0;
      type_cast_2512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2512_inst_req_1;
      type_cast_2512_inst_ack_1<= rack(0);
      type_cast_2512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2528_inst_req_0;
      type_cast_2528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2528_inst_req_1;
      type_cast_2528_inst_ack_1<= rack(0);
      type_cast_2528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2545_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2545_inst_req_0;
      type_cast_2545_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2545_inst_req_1;
      type_cast_2545_inst_ack_1<= rack(0);
      type_cast_2545_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2545_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2496,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2545_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2552_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2552_inst_req_0;
      type_cast_2552_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2552_inst_req_1;
      type_cast_2552_inst_ack_1<= rack(0);
      type_cast_2552_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2552_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2552_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2554_inst_req_0;
      type_cast_2554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2554_inst_req_1;
      type_cast_2554_inst_ack_1<= rack(0);
      type_cast_2554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2554_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2558_inst_req_0;
      type_cast_2558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2558_inst_req_1;
      type_cast_2558_inst_ack_1<= rack(0);
      type_cast_2558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2558_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2560_inst_req_0;
      type_cast_2560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2560_inst_req_1;
      type_cast_2560_inst_ack_1<= rack(0);
      type_cast_2560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2560_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2439_index_1_rename
    process(R_idxprom_2438_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2438_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2438_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2439_index_1_resize
    process(idxprom_2434) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2434;
      ov := iv(13 downto 0);
      R_idxprom_2438_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2439_root_address_inst
    process(array_obj_ref_2439_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2439_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2439_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2462_index_1_rename
    process(R_idxprom86_2461_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2461_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2461_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2462_index_1_resize
    process(idxprom86_2457) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2457;
      ov := iv(13 downto 0);
      R_idxprom86_2461_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2462_root_address_inst
    process(array_obj_ref_2462_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2462_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2462_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2444_addr_0
    process(ptr_deref_2444_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2444_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2444_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2444_base_resize
    process(arrayidx82_2441) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2441;
      ov := iv(13 downto 0);
      ptr_deref_2444_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2444_gather_scatter
    process(ptr_deref_2444_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2444_data_0;
      ov(63 downto 0) := iv;
      tmp83_2445 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2444_root_address_inst
    process(ptr_deref_2444_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2444_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2444_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2466_addr_0
    process(ptr_deref_2466_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2466_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2466_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2466_base_resize
    process(arrayidx87_2464) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2464;
      ov := iv(13 downto 0);
      ptr_deref_2466_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2466_gather_scatter
    process(tmp83_2445) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2445;
      ov(63 downto 0) := iv;
      ptr_deref_2466_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2466_root_address_inst
    process(ptr_deref_2466_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2466_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2466_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2484_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2483;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2484_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2484_branch_req_0,
          ack0 => if_stmt_2484_branch_ack_0,
          ack1 => if_stmt_2484_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2535_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2534;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2535_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2535_branch_req_0,
          ack0 => if_stmt_2535_branch_ack_0,
          ack1 => if_stmt_2535_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2281_inst
    process(call7_2223) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2223, type_cast_2280_wire_constant, tmp_var);
      add45_2282 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2292_inst
    process(call9_2226) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2226, type_cast_2291_wire_constant, tmp_var);
      add58_2293 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2381_inst
    process(sub_2287, mul_2377) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2287, mul_2377, tmp_var);
      sub48_2382 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2391_inst
    process(sub61_2298, mul54_2387) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2298, mul54_2387, tmp_var);
      sub62_2392 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2495_inst
    process(input_dim2x_x1_2341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2341, type_cast_2494_wire_constant, tmp_var);
      add98_2496 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2503_inst
    process(input_dim1x_x1_2348) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2348, type_cast_2502_wire_constant, tmp_var);
      inc_2504 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2517_inst
    process(inc110_2513, input_dim0x_x2_2355) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2513, input_dim0x_x2_2355, tmp_var);
      inc110x_xinput_dim0x_x2_2518 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2330_inst
    process(shr116137_2320, shr120138_2326) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2320, shr120138_2326, tmp_var);
      add121_2331 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2371_inst
    process(add_2260, tmp1_2367) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2260, tmp1_2367, tmp_var);
      add_src_0x_x0_2372 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2477_inst
    process(conv90_2472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2472, type_cast_2476_wire_constant, tmp_var);
      add91_2478 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2566_inst
    process(indvar_2334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2334, type_cast_2565_wire_constant, tmp_var);
      indvarx_xnext_2567 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2413_inst
    process(mul76_2409, conv70_2400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2409, conv70_2400, tmp_var);
      add77_2414 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2423_inst
    process(mul78_2419, conv65_2396) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2419, conv65_2396, tmp_var);
      add79_2424 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2456_inst
    process(shr85_2451) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2451, type_cast_2455_wire_constant, tmp_var);
      idxprom86_2457 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2508_inst
    process(inc_2504, call1_2214) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2504, call1_2214, tmp_var);
      cmp106_2509 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2533_inst
    process(conv112_2529, add121_2331) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2529, add121_2331, tmp_var);
      cmp122_2534 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2275_inst
    process(call_2211) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2211, type_cast_2274_wire_constant, tmp_var);
      shr136_2276 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2319_inst
    process(conv115_2314) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2314, type_cast_2318_wire_constant, tmp_var);
      shr116137_2320 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2325_inst
    process(conv115_2314) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2314, type_cast_2324_wire_constant, tmp_var);
      shr120138_2326 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2429_inst
    process(add_src_0x_x0_2372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2372, type_cast_2428_wire_constant, tmp_var);
      shr81_2430 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2450_inst
    process(add79_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2424, type_cast_2449_wire_constant, tmp_var);
      shr85_2451 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2376_inst
    process(input_dim0x_x2_2355, call13_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2355, call13_2232, tmp_var);
      mul_2377 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2386_inst
    process(input_dim1x_x1_2348, call13_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2348, call13_2232, tmp_var);
      mul54_2387 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2366_inst
    process(indvar_2334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2334, type_cast_2365_wire_constant, tmp_var);
      tmp1_2367 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2408_inst
    process(conv75_2404, conv73_2306) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2404, conv73_2306, tmp_var);
      mul76_2409 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2418_inst
    process(add77_2414, conv68_2302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2414, conv68_2302, tmp_var);
      mul78_2419 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2259_inst
    process(shl_2248, conv17_2255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2248, conv17_2255, tmp_var);
      add_2260 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2247_inst
    process(conv_2242) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2242, type_cast_2246_wire_constant, tmp_var);
      shl_2248 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2286_inst
    process(add45_2282, call14_2235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2282, call14_2235, tmp_var);
      sub_2287 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2297_inst
    process(add58_2293, call14_2235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2293, call14_2235, tmp_var);
      sub61_2298 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2482_inst
    process(add91_2478, conv94_2310) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2478, conv94_2310, tmp_var);
      cmp_2483 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2439_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2438_scaled;
      array_obj_ref_2439_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2439_index_offset_req_0;
      array_obj_ref_2439_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2439_index_offset_req_1;
      array_obj_ref_2439_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2462_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2461_scaled;
      array_obj_ref_2462_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2462_index_offset_req_0;
      array_obj_ref_2462_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2462_index_offset_req_1;
      array_obj_ref_2462_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2444_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2444_load_0_req_0;
      ptr_deref_2444_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2444_load_0_req_1;
      ptr_deref_2444_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2444_word_address_0;
      ptr_deref_2444_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2466_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2466_store_0_req_0;
      ptr_deref_2466_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2466_store_0_req_1;
      ptr_deref_2466_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2466_word_address_0;
      data_in <= ptr_deref_2466_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2250_inst RPIPE_Block2_start_2262_inst RPIPE_Block2_start_2265_inst RPIPE_Block2_start_2268_inst RPIPE_Block2_start_2237_inst RPIPE_Block2_start_2234_inst RPIPE_Block2_start_2231_inst RPIPE_Block2_start_2228_inst RPIPE_Block2_start_2225_inst RPIPE_Block2_start_2222_inst RPIPE_Block2_start_2219_inst RPIPE_Block2_start_2216_inst RPIPE_Block2_start_2213_inst RPIPE_Block2_start_2210_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2250_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2262_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2265_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2268_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2237_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2234_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2231_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2228_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2225_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2222_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2219_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2216_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2213_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2210_inst_req_0;
      RPIPE_Block2_start_2250_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2262_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2265_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2268_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2237_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2234_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2231_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2228_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2225_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2222_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2219_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2216_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2213_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2210_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2250_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2262_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2265_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2268_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2237_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2234_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2231_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2228_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2225_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2222_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2219_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2216_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2213_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2210_inst_req_1;
      RPIPE_Block2_start_2250_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2262_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2265_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2268_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2237_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2234_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2231_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2228_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2225_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2222_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2219_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2216_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2213_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2210_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call16_2251 <= data_out(223 downto 208);
      call18_2263 <= data_out(207 downto 192);
      call20_2266 <= data_out(191 downto 176);
      call22_2269 <= data_out(175 downto 160);
      call15_2238 <= data_out(159 downto 144);
      call14_2235 <= data_out(143 downto 128);
      call13_2232 <= data_out(127 downto 112);
      call11_2229 <= data_out(111 downto 96);
      call9_2226 <= data_out(95 downto 80);
      call7_2223 <= data_out(79 downto 64);
      call5_2220 <= data_out(63 downto 48);
      call3_2217 <= data_out(47 downto 32);
      call1_2214 <= data_out(31 downto 16);
      call_2211 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2571_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2571_inst_req_0;
      WPIPE_Block2_done_2571_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2571_inst_req_1;
      WPIPE_Block2_done_2571_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2573_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6773_start: Boolean;
  signal convTransposeD_CP_6773_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2640_inst_ack_1 : boolean;
  signal type_cast_2692_inst_ack_0 : boolean;
  signal type_cast_2692_inst_req_0 : boolean;
  signal type_cast_2795_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2622_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2637_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2640_inst_req_1 : boolean;
  signal type_cast_2761_inst_ack_0 : boolean;
  signal type_cast_2761_inst_ack_1 : boolean;
  signal array_obj_ref_2801_index_offset_ack_0 : boolean;
  signal RPIPE_Block3_start_2637_inst_req_0 : boolean;
  signal type_cast_2761_inst_req_1 : boolean;
  signal type_cast_2688_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2637_inst_ack_0 : boolean;
  signal addr_of_2802_final_reg_ack_1 : boolean;
  signal type_cast_2765_inst_req_0 : boolean;
  signal type_cast_2757_inst_ack_1 : boolean;
  signal type_cast_2626_inst_req_1 : boolean;
  signal array_obj_ref_2801_index_offset_req_0 : boolean;
  signal addr_of_2802_final_reg_req_1 : boolean;
  signal RPIPE_Block3_start_2634_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2622_inst_req_1 : boolean;
  signal type_cast_2795_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2640_inst_req_0 : boolean;
  signal type_cast_2626_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2634_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2640_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2634_inst_req_1 : boolean;
  signal type_cast_2688_inst_req_0 : boolean;
  signal type_cast_2757_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2634_inst_ack_1 : boolean;
  signal array_obj_ref_2801_index_offset_req_1 : boolean;
  signal type_cast_2795_inst_req_1 : boolean;
  signal type_cast_2688_inst_ack_0 : boolean;
  signal type_cast_2692_inst_req_1 : boolean;
  signal type_cast_2684_inst_req_0 : boolean;
  signal type_cast_2692_inst_ack_1 : boolean;
  signal array_obj_ref_2801_index_offset_ack_1 : boolean;
  signal type_cast_2757_inst_req_0 : boolean;
  signal type_cast_2765_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2622_inst_ack_1 : boolean;
  signal type_cast_2684_inst_req_1 : boolean;
  signal type_cast_2765_inst_req_1 : boolean;
  signal type_cast_2757_inst_ack_0 : boolean;
  signal type_cast_2626_inst_req_0 : boolean;
  signal type_cast_2688_inst_req_1 : boolean;
  signal type_cast_2765_inst_ack_1 : boolean;
  signal addr_of_2802_final_reg_req_0 : boolean;
  signal type_cast_2626_inst_ack_0 : boolean;
  signal type_cast_2613_inst_req_1 : boolean;
  signal addr_of_2802_final_reg_ack_0 : boolean;
  signal type_cast_2684_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2622_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2637_inst_ack_1 : boolean;
  signal type_cast_2613_inst_ack_1 : boolean;
  signal type_cast_2684_inst_ack_0 : boolean;
  signal type_cast_2795_inst_ack_1 : boolean;
  signal type_cast_2761_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2582_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2582_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2582_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2582_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2585_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2585_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2585_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2585_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2591_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2591_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2591_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2591_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2594_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2594_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2594_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2594_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2597_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2597_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2597_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2597_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2600_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2600_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2600_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2600_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2603_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2603_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2603_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2603_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2609_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2609_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2609_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2609_inst_ack_1 : boolean;
  signal type_cast_2613_inst_req_0 : boolean;
  signal type_cast_2613_inst_ack_0 : boolean;
  signal ptr_deref_2806_load_0_req_0 : boolean;
  signal ptr_deref_2806_load_0_ack_0 : boolean;
  signal ptr_deref_2806_load_0_req_1 : boolean;
  signal ptr_deref_2806_load_0_ack_1 : boolean;
  signal array_obj_ref_2824_index_offset_req_0 : boolean;
  signal array_obj_ref_2824_index_offset_ack_0 : boolean;
  signal array_obj_ref_2824_index_offset_req_1 : boolean;
  signal array_obj_ref_2824_index_offset_ack_1 : boolean;
  signal addr_of_2825_final_reg_req_0 : boolean;
  signal addr_of_2825_final_reg_ack_0 : boolean;
  signal addr_of_2825_final_reg_req_1 : boolean;
  signal addr_of_2825_final_reg_ack_1 : boolean;
  signal ptr_deref_2828_store_0_req_0 : boolean;
  signal ptr_deref_2828_store_0_ack_0 : boolean;
  signal ptr_deref_2828_store_0_req_1 : boolean;
  signal ptr_deref_2828_store_0_ack_1 : boolean;
  signal type_cast_2833_inst_req_0 : boolean;
  signal type_cast_2833_inst_ack_0 : boolean;
  signal type_cast_2833_inst_req_1 : boolean;
  signal type_cast_2833_inst_ack_1 : boolean;
  signal if_stmt_2846_branch_req_0 : boolean;
  signal if_stmt_2846_branch_ack_1 : boolean;
  signal if_stmt_2846_branch_ack_0 : boolean;
  signal type_cast_2874_inst_req_0 : boolean;
  signal type_cast_2874_inst_ack_0 : boolean;
  signal type_cast_2874_inst_req_1 : boolean;
  signal type_cast_2874_inst_ack_1 : boolean;
  signal if_stmt_2893_branch_req_0 : boolean;
  signal if_stmt_2893_branch_ack_1 : boolean;
  signal if_stmt_2893_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2929_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2929_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2929_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2929_inst_ack_1 : boolean;
  signal phi_stmt_2696_req_0 : boolean;
  signal phi_stmt_2703_req_0 : boolean;
  signal phi_stmt_2710_req_0 : boolean;
  signal type_cast_2720_inst_req_0 : boolean;
  signal type_cast_2720_inst_ack_0 : boolean;
  signal type_cast_2720_inst_req_1 : boolean;
  signal type_cast_2720_inst_ack_1 : boolean;
  signal phi_stmt_2717_req_0 : boolean;
  signal type_cast_2702_inst_req_0 : boolean;
  signal type_cast_2702_inst_ack_0 : boolean;
  signal type_cast_2702_inst_req_1 : boolean;
  signal type_cast_2702_inst_ack_1 : boolean;
  signal phi_stmt_2696_req_1 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal phi_stmt_2703_req_1 : boolean;
  signal type_cast_2716_inst_req_0 : boolean;
  signal type_cast_2716_inst_ack_0 : boolean;
  signal type_cast_2716_inst_req_1 : boolean;
  signal type_cast_2716_inst_ack_1 : boolean;
  signal phi_stmt_2710_req_1 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal phi_stmt_2717_req_1 : boolean;
  signal phi_stmt_2696_ack_0 : boolean;
  signal phi_stmt_2703_ack_0 : boolean;
  signal phi_stmt_2710_ack_0 : boolean;
  signal phi_stmt_2717_ack_0 : boolean;
  signal phi_stmt_2900_req_1 : boolean;
  signal type_cast_2912_inst_req_0 : boolean;
  signal type_cast_2912_inst_ack_0 : boolean;
  signal type_cast_2912_inst_req_1 : boolean;
  signal type_cast_2912_inst_ack_1 : boolean;
  signal phi_stmt_2907_req_1 : boolean;
  signal type_cast_2918_inst_req_0 : boolean;
  signal type_cast_2918_inst_ack_0 : boolean;
  signal type_cast_2918_inst_req_1 : boolean;
  signal type_cast_2918_inst_ack_1 : boolean;
  signal phi_stmt_2913_req_1 : boolean;
  signal type_cast_2903_inst_req_0 : boolean;
  signal type_cast_2903_inst_ack_0 : boolean;
  signal type_cast_2903_inst_req_1 : boolean;
  signal type_cast_2903_inst_ack_1 : boolean;
  signal phi_stmt_2900_req_0 : boolean;
  signal type_cast_2910_inst_req_0 : boolean;
  signal type_cast_2910_inst_ack_0 : boolean;
  signal type_cast_2910_inst_req_1 : boolean;
  signal type_cast_2910_inst_ack_1 : boolean;
  signal phi_stmt_2907_req_0 : boolean;
  signal type_cast_2916_inst_req_0 : boolean;
  signal type_cast_2916_inst_ack_0 : boolean;
  signal type_cast_2916_inst_req_1 : boolean;
  signal type_cast_2916_inst_ack_1 : boolean;
  signal phi_stmt_2913_req_0 : boolean;
  signal phi_stmt_2900_ack_0 : boolean;
  signal phi_stmt_2907_ack_0 : boolean;
  signal phi_stmt_2913_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6773_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6773: Block -- control-path 
    signal convTransposeD_CP_6773_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6773_elements(0) <= convTransposeD_CP_6773_start;
    convTransposeD_CP_6773_symbol <= convTransposeD_CP_6773_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2580/$entry
      -- CP-element group 0: 	 branch_block_stmt_2580/branch_block_stmt_2580__entry__
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641__entry__
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/$entry
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_update_start_
      -- 
    cr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => type_cast_2626_inst_req_1); -- 
    cr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => type_cast_2613_inst_req_1); -- 
    rr_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => RPIPE_Block3_start_2582_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2580/merge_stmt_2899__exit__
      -- CP-element group 1: 	 branch_block_stmt_2580/assign_stmt_2925__entry__
      -- CP-element group 1: 	 branch_block_stmt_2580/assign_stmt_2925__exit__
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2580/assign_stmt_2925/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/assign_stmt_2925/$exit
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Update/cr
      -- 
    rr_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2702_inst_req_0); -- 
    cr_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2702_inst_req_1); -- 
    rr_7517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2709_inst_req_0); -- 
    cr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2709_inst_req_1); -- 
    rr_7540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2716_inst_req_0); -- 
    cr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2716_inst_req_1); -- 
    rr_7563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2722_inst_req_0); -- 
    cr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2722_inst_req_1); -- 
    convTransposeD_CP_6773_elements(1) <= convTransposeD_CP_6773_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Update/cr
      -- 
    ra_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2582_inst_ack_0, ack => convTransposeD_CP_6773_elements(2)); -- 
    cr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(2), ack => RPIPE_Block3_start_2582_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2582_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Sample/rr
      -- 
    ca_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2582_inst_ack_1, ack => convTransposeD_CP_6773_elements(3)); -- 
    rr_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(3), ack => RPIPE_Block3_start_2585_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Update/cr
      -- 
    ra_6836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2585_inst_ack_0, ack => convTransposeD_CP_6773_elements(4)); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(4), ack => RPIPE_Block3_start_2585_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2585_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Sample/rr
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2585_inst_ack_1, ack => convTransposeD_CP_6773_elements(5)); -- 
    rr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(5), ack => RPIPE_Block3_start_2588_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Update/cr
      -- 
    ra_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_0, ack => convTransposeD_CP_6773_elements(6)); -- 
    cr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(6), ack => RPIPE_Block3_start_2588_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2588_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Sample/rr
      -- 
    ca_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_1, ack => convTransposeD_CP_6773_elements(7)); -- 
    rr_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(7), ack => RPIPE_Block3_start_2591_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Update/cr
      -- 
    ra_6864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2591_inst_ack_0, ack => convTransposeD_CP_6773_elements(8)); -- 
    cr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(8), ack => RPIPE_Block3_start_2591_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2591_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Sample/rr
      -- 
    ca_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2591_inst_ack_1, ack => convTransposeD_CP_6773_elements(9)); -- 
    rr_6877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(9), ack => RPIPE_Block3_start_2594_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Update/cr
      -- 
    ra_6878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2594_inst_ack_0, ack => convTransposeD_CP_6773_elements(10)); -- 
    cr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(10), ack => RPIPE_Block3_start_2594_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2594_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Sample/rr
      -- 
    ca_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2594_inst_ack_1, ack => convTransposeD_CP_6773_elements(11)); -- 
    rr_6891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(11), ack => RPIPE_Block3_start_2597_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Update/cr
      -- 
    ra_6892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2597_inst_ack_0, ack => convTransposeD_CP_6773_elements(12)); -- 
    cr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(12), ack => RPIPE_Block3_start_2597_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2597_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Sample/rr
      -- 
    ca_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2597_inst_ack_1, ack => convTransposeD_CP_6773_elements(13)); -- 
    rr_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(13), ack => RPIPE_Block3_start_2600_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Update/cr
      -- 
    ra_6906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2600_inst_ack_0, ack => convTransposeD_CP_6773_elements(14)); -- 
    cr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(14), ack => RPIPE_Block3_start_2600_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2600_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Sample/rr
      -- 
    ca_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2600_inst_ack_1, ack => convTransposeD_CP_6773_elements(15)); -- 
    rr_6919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(15), ack => RPIPE_Block3_start_2603_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Update/cr
      -- 
    ra_6920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2603_inst_ack_0, ack => convTransposeD_CP_6773_elements(16)); -- 
    cr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(16), ack => RPIPE_Block3_start_2603_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2603_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Sample/rr
      -- 
    ca_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2603_inst_ack_1, ack => convTransposeD_CP_6773_elements(17)); -- 
    rr_6933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(17), ack => RPIPE_Block3_start_2606_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Update/cr
      -- 
    ra_6934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_0, ack => convTransposeD_CP_6773_elements(18)); -- 
    cr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(18), ack => RPIPE_Block3_start_2606_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2606_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Sample/rr
      -- 
    ca_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_1, ack => convTransposeD_CP_6773_elements(19)); -- 
    rr_6947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(19), ack => RPIPE_Block3_start_2609_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Update/cr
      -- 
    ra_6948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2609_inst_ack_0, ack => convTransposeD_CP_6773_elements(20)); -- 
    cr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(20), ack => RPIPE_Block3_start_2609_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2609_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Sample/rr
      -- 
    ca_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2609_inst_ack_1, ack => convTransposeD_CP_6773_elements(21)); -- 
    rr_6961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(21), ack => type_cast_2613_inst_req_0); -- 
    rr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(21), ack => RPIPE_Block3_start_2622_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Sample/ra
      -- 
    ra_6962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_0, ack => convTransposeD_CP_6773_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2613_update_completed_
      -- 
    ca_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2613_inst_ack_1, ack => convTransposeD_CP_6773_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Update/$entry
      -- 
    ra_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2622_inst_ack_0, ack => convTransposeD_CP_6773_elements(24)); -- 
    cr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(24), ack => RPIPE_Block3_start_2622_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2622_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Sample/rr
      -- 
    ca_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2622_inst_ack_1, ack => convTransposeD_CP_6773_elements(25)); -- 
    rr_6989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(25), ack => type_cast_2626_inst_req_0); -- 
    rr_7003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(25), ack => RPIPE_Block3_start_2634_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Sample/ra
      -- 
    ra_6990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2626_inst_ack_0, ack => convTransposeD_CP_6773_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/type_cast_2626_Update/ca
      -- 
    ca_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2626_inst_ack_1, ack => convTransposeD_CP_6773_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_update_start_
      -- 
    ra_7004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2634_inst_ack_0, ack => convTransposeD_CP_6773_elements(28)); -- 
    cr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(28), ack => RPIPE_Block3_start_2634_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2634_Update/ca
      -- 
    ca_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2634_inst_ack_1, ack => convTransposeD_CP_6773_elements(29)); -- 
    rr_7017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(29), ack => RPIPE_Block3_start_2637_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Update/$entry
      -- 
    ra_7018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2637_inst_ack_0, ack => convTransposeD_CP_6773_elements(30)); -- 
    cr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(30), ack => RPIPE_Block3_start_2637_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2637_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_sample_start_
      -- 
    ca_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2637_inst_ack_1, ack => convTransposeD_CP_6773_elements(31)); -- 
    rr_7031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(31), ack => RPIPE_Block3_start_2640_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Update/$entry
      -- 
    ra_7032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2640_inst_ack_0, ack => convTransposeD_CP_6773_elements(32)); -- 
    cr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(32), ack => RPIPE_Block3_start_2640_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/RPIPE_Block3_start_2640_Update/$exit
      -- 
    ca_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2640_inst_ack_1, ack => convTransposeD_CP_6773_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641__exit__
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693__entry__
      -- CP-element group 34: 	 branch_block_stmt_2580/assign_stmt_2583_to_assign_stmt_2641/$exit
      -- 
    rr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2692_inst_req_0); -- 
    rr_7062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2688_inst_req_0); -- 
    cr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2692_inst_req_1); -- 
    rr_7048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2684_inst_req_0); -- 
    cr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2684_inst_req_1); -- 
    cr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2688_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(23) & convTransposeD_CP_6773_elements(27) & convTransposeD_CP_6773_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Sample/ra
      -- 
    ra_7049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_0, ack => convTransposeD_CP_6773_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2684_Update/ca
      -- 
    ca_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_1, ack => convTransposeD_CP_6773_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Sample/ra
      -- 
    ra_7063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2688_inst_ack_0, ack => convTransposeD_CP_6773_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2688_Update/$exit
      -- 
    ca_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2688_inst_ack_1, ack => convTransposeD_CP_6773_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_sample_completed_
      -- 
    ra_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_0, ack => convTransposeD_CP_6773_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/type_cast_2692_Update/ca
      -- 
    ca_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_1, ack => convTransposeD_CP_6773_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693/$exit
      -- CP-element group 41: 	 branch_block_stmt_2580/assign_stmt_2648_to_assign_stmt_2693__exit__
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Update/cr
      -- 
    rr_7468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(41), ack => type_cast_2720_inst_req_0); -- 
    cr_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(41), ack => type_cast_2720_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(36) & convTransposeD_CP_6773_elements(38) & convTransposeD_CP_6773_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_sample_completed_
      -- 
    ra_7094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2757_inst_ack_0, ack => convTransposeD_CP_6773_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Update/$exit
      -- 
    ca_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2757_inst_ack_1, ack => convTransposeD_CP_6773_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Sample/$exit
      -- 
    ra_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2761_inst_ack_0, ack => convTransposeD_CP_6773_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Update/$exit
      -- 
    ca_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2761_inst_ack_1, ack => convTransposeD_CP_6773_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Sample/ra
      -- 
    ra_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2765_inst_ack_0, ack => convTransposeD_CP_6773_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Update/$exit
      -- 
    ca_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2765_inst_ack_1, ack => convTransposeD_CP_6773_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_sample_completed_
      -- 
    ra_7136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_0, ack => convTransposeD_CP_6773_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Update/ca
      -- 
    ca_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2795_inst_ack_1, ack => convTransposeD_CP_6773_elements(49)); -- 
    req_7166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(49), ack => array_obj_ref_2801_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_sample_complete
      -- 
    ack_7167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2801_index_offset_ack_0, ack => convTransposeD_CP_6773_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_request/req
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_sample_start_
      -- 
    ack_7172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2801_index_offset_ack_1, ack => convTransposeD_CP_6773_elements(51)); -- 
    req_7181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(51), ack => addr_of_2802_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_request/ack
      -- CP-element group 52: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_request/$exit
      -- 
    ack_7182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2802_final_reg_ack_0, ack => convTransposeD_CP_6773_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/word_0/rr
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2802_final_reg_ack_1, ack => convTransposeD_CP_6773_elements(53)); -- 
    rr_7220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(53), ack => ptr_deref_2806_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Sample/word_access_start/word_0/ra
      -- 
    ra_7221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2806_load_0_ack_0, ack => convTransposeD_CP_6773_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/ptr_deref_2806_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/ptr_deref_2806_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/ptr_deref_2806_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/ptr_deref_2806_Merge/merge_ack
      -- 
    ca_7232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2806_load_0_ack_1, ack => convTransposeD_CP_6773_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Sample/req
      -- 
    req_7262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(56), ack => array_obj_ref_2824_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(43) & convTransposeD_CP_6773_elements(45) & convTransposeD_CP_6773_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Sample/ack
      -- 
    ack_7263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2824_index_offset_ack_0, ack => convTransposeD_CP_6773_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_request/req
      -- 
    ack_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2824_index_offset_ack_1, ack => convTransposeD_CP_6773_elements(58)); -- 
    req_7277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(58), ack => addr_of_2825_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_request/ack
      -- 
    ack_7278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2825_final_reg_ack_0, ack => convTransposeD_CP_6773_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_word_addrgen/root_register_ack
      -- 
    ack_7283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2825_final_reg_ack_1, ack => convTransposeD_CP_6773_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/ptr_deref_2828_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/ptr_deref_2828_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/ptr_deref_2828_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/ptr_deref_2828_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/word_0/rr
      -- 
    rr_7321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(61), ack => ptr_deref_2828_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(55) & convTransposeD_CP_6773_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Sample/word_access_start/word_0/ra
      -- 
    ra_7322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2828_store_0_ack_0, ack => convTransposeD_CP_6773_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/word_0/ca
      -- 
    ca_7333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2828_store_0_ack_1, ack => convTransposeD_CP_6773_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Sample/ra
      -- 
    ra_7342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2833_inst_ack_0, ack => convTransposeD_CP_6773_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Update/ca
      -- 
    ca_7347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2833_inst_ack_1, ack => convTransposeD_CP_6773_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2580/R_cmp_2847_place
      -- CP-element group 66: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/$exit
      -- CP-element group 66: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845__exit__
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846__entry__
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2580/if_stmt_2846_else_link/$entry
      -- 
    branch_req_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(66), ack => if_stmt_2846_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(50) & convTransposeD_CP_6773_elements(57) & convTransposeD_CP_6773_elements(63) & convTransposeD_CP_6773_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2580/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2580/merge_stmt_2852__exit__
      -- CP-element group 67: 	 branch_block_stmt_2580/assign_stmt_2858__entry__
      -- CP-element group 67: 	 branch_block_stmt_2580/assign_stmt_2858__exit__
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2580/if_stmt_2846_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2580/if_stmt_2846_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2580/assign_stmt_2858/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/assign_stmt_2858/$exit
      -- CP-element group 67: 	 branch_block_stmt_2580/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2580/merge_stmt_2852_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2580/merge_stmt_2852_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/merge_stmt_2852_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2580/merge_stmt_2852_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2846_branch_ack_1, ack => convTransposeD_CP_6773_elements(67)); -- 
    rr_7678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2903_inst_req_0); -- 
    cr_7683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2903_inst_req_1); -- 
    rr_7701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2910_inst_req_0); -- 
    cr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2910_inst_req_1); -- 
    rr_7724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2916_inst_req_0); -- 
    cr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2916_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2580/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2580/merge_stmt_2860__exit__
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892__entry__
      -- CP-element group 68: 	 branch_block_stmt_2580/if_stmt_2846_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2580/if_stmt_2846_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/$entry
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2580/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2580/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2580/merge_stmt_2860_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2580/merge_stmt_2860_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2580/merge_stmt_2860_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2580/merge_stmt_2860_PhiAck/dummy
      -- 
    else_choice_transition_7364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2846_branch_ack_0, ack => convTransposeD_CP_6773_elements(68)); -- 
    rr_7380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(68), ack => type_cast_2874_inst_req_0); -- 
    cr_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(68), ack => type_cast_2874_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Sample/ra
      -- 
    ra_7381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_0, ack => convTransposeD_CP_6773_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892__exit__
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893__entry__
      -- CP-element group 70: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/$exit
      -- CP-element group 70: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2580/assign_stmt_2866_to_assign_stmt_2892/type_cast_2874_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2580/R_cmp121_2894_place
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2580/if_stmt_2893_else_link/$entry
      -- 
    ca_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2874_inst_ack_1, ack => convTransposeD_CP_6773_elements(70)); -- 
    branch_req_7394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(70), ack => if_stmt_2893_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2580/merge_stmt_2927__exit__
      -- CP-element group 71: 	 branch_block_stmt_2580/assign_stmt_2932__entry__
      -- CP-element group 71: 	 branch_block_stmt_2580/if_stmt_2893_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2580/if_stmt_2893_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2580/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2580/assign_stmt_2932/$entry
      -- CP-element group 71: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2580/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2580/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2580/merge_stmt_2927_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2580/merge_stmt_2927_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2580/merge_stmt_2927_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2580/merge_stmt_2927_PhiAck/dummy
      -- 
    if_choice_transition_7399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2893_branch_ack_1, ack => convTransposeD_CP_6773_elements(71)); -- 
    req_7419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(71), ack => WPIPE_Block3_done_2929_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2580/if_stmt_2893_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2580/if_stmt_2893_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2893_branch_ack_0, ack => convTransposeD_CP_6773_elements(72)); -- 
    rr_7629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2912_inst_req_0); -- 
    cr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2912_inst_req_1); -- 
    rr_7652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2918_inst_req_0); -- 
    cr_7657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2918_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Update/req
      -- 
    ack_7420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2929_inst_ack_0, ack => convTransposeD_CP_6773_elements(73)); -- 
    req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(73), ack => WPIPE_Block3_done_2929_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2580/$exit
      -- CP-element group 74: 	 branch_block_stmt_2580/branch_block_stmt_2580__exit__
      -- CP-element group 74: 	 branch_block_stmt_2580/assign_stmt_2932__exit__
      -- CP-element group 74: 	 branch_block_stmt_2580/return__
      -- CP-element group 74: 	 branch_block_stmt_2580/merge_stmt_2934__exit__
      -- CP-element group 74: 	 branch_block_stmt_2580/assign_stmt_2932/$exit
      -- CP-element group 74: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2580/assign_stmt_2932/WPIPE_Block3_done_2929_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2580/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2580/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2580/merge_stmt_2934_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2580/merge_stmt_2934_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2580/merge_stmt_2934_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2580/merge_stmt_2934_PhiAck/dummy
      -- 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2929_inst_ack_1, ack => convTransposeD_CP_6773_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/$exit
      -- CP-element group 75: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2700_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_req
      -- 
    phi_stmt_2696_req_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2696_req_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(75), ack => phi_stmt_2696_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/$exit
      -- CP-element group 76: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2707_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_req
      -- 
    phi_stmt_2703_req_7444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2703_req_7444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(76), ack => phi_stmt_2703_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/$exit
      -- CP-element group 77: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2714_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_req
      -- 
    phi_stmt_2710_req_7452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2710_req_7452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(77), ack => phi_stmt_2710_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Sample/ra
      -- 
    ra_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2720_inst_ack_0, ack => convTransposeD_CP_6773_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/Update/ca
      -- 
    ca_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2720_inst_ack_1, ack => convTransposeD_CP_6773_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/$exit
      -- CP-element group 80: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/$exit
      -- CP-element group 80: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2720/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_req
      -- 
    phi_stmt_2717_req_7475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2717_req_7475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(80), ack => phi_stmt_2717_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(78) & convTransposeD_CP_6773_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2580/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(75) & convTransposeD_CP_6773_elements(76) & convTransposeD_CP_6773_elements(77) & convTransposeD_CP_6773_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Sample/ra
      -- 
    ra_7495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2702_inst_ack_0, ack => convTransposeD_CP_6773_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/Update/ca
      -- 
    ca_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2702_inst_ack_1, ack => convTransposeD_CP_6773_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/$exit
      -- CP-element group 84: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/$exit
      -- CP-element group 84: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_sources/type_cast_2702/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2696/phi_stmt_2696_req
      -- 
    phi_stmt_2696_req_7501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2696_req_7501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(84), ack => phi_stmt_2696_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(82) & convTransposeD_CP_6773_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Sample/ra
      -- 
    ra_7518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => convTransposeD_CP_6773_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/Update/ca
      -- 
    ca_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => convTransposeD_CP_6773_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/$exit
      -- CP-element group 87: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/$exit
      -- CP-element group 87: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_sources/type_cast_2709/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2703/phi_stmt_2703_req
      -- 
    phi_stmt_2703_req_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2703_req_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(87), ack => phi_stmt_2703_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(85) & convTransposeD_CP_6773_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Sample/ra
      -- 
    ra_7541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2716_inst_ack_0, ack => convTransposeD_CP_6773_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/Update/ca
      -- 
    ca_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2716_inst_ack_1, ack => convTransposeD_CP_6773_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/$exit
      -- CP-element group 90: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/$exit
      -- CP-element group 90: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_sources/type_cast_2716/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2710/phi_stmt_2710_req
      -- 
    phi_stmt_2710_req_7547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2710_req_7547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(90), ack => phi_stmt_2710_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(88) & convTransposeD_CP_6773_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Sample/ra
      -- 
    ra_7564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeD_CP_6773_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/Update/ca
      -- 
    ca_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeD_CP_6773_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/$exit
      -- CP-element group 93: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/$exit
      -- CP-element group 93: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_sources/type_cast_2722/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2717/phi_stmt_2717_req
      -- 
    phi_stmt_2717_req_7570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2717_req_7570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(93), ack => phi_stmt_2717_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(91) & convTransposeD_CP_6773_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2580/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(84) & convTransposeD_CP_6773_elements(87) & convTransposeD_CP_6773_elements(90) & convTransposeD_CP_6773_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2580/merge_stmt_2695_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/$entry
      -- 
    convTransposeD_CP_6773_elements(95) <= OrReduce(convTransposeD_CP_6773_elements(81) & convTransposeD_CP_6773_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/phi_stmt_2696_ack
      -- 
    phi_stmt_2696_ack_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2696_ack_0, ack => convTransposeD_CP_6773_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/phi_stmt_2703_ack
      -- 
    phi_stmt_2703_ack_7576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2703_ack_0, ack => convTransposeD_CP_6773_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/phi_stmt_2710_ack
      -- 
    phi_stmt_2710_ack_7577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2710_ack_0, ack => convTransposeD_CP_6773_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/phi_stmt_2717_ack
      -- 
    phi_stmt_2717_ack_7578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2717_ack_0, ack => convTransposeD_CP_6773_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2765_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2802_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2801_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2757_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2761_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2580/merge_stmt_2695__exit__
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845__entry__
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2795_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2806_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/array_obj_ref_2824_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/addr_of_2825_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/ptr_deref_2828_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2580/assign_stmt_2729_to_assign_stmt_2845/type_cast_2833_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2580/merge_stmt_2695_PhiAck/$exit
      -- 
    rr_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2795_inst_req_0); -- 
    cr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2761_inst_req_1); -- 
    rr_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2765_inst_req_0); -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => addr_of_2802_final_reg_req_1); -- 
    cr_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2757_inst_req_1); -- 
    req_7171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => array_obj_ref_2801_index_offset_req_1); -- 
    cr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2795_inst_req_1); -- 
    rr_7093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2757_inst_req_0); -- 
    cr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2765_inst_req_1); -- 
    rr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2761_inst_req_0); -- 
    cr_7231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => ptr_deref_2806_load_0_req_1); -- 
    req_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => array_obj_ref_2824_index_offset_req_1); -- 
    req_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => addr_of_2825_final_reg_req_1); -- 
    cr_7332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => ptr_deref_2828_store_0_req_1); -- 
    rr_7341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2833_inst_req_0); -- 
    cr_7346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2833_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(96) & convTransposeD_CP_6773_elements(97) & convTransposeD_CP_6773_elements(98) & convTransposeD_CP_6773_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/$exit
      -- CP-element group 101: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2906_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_req
      -- 
    phi_stmt_2900_req_7613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2900_req_7613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(101), ack => phi_stmt_2900_req_1); -- 
    -- Element group convTransposeD_CP_6773_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(72), ack => convTransposeD_CP_6773_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Sample/ra
      -- 
    ra_7630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2912_inst_ack_0, ack => convTransposeD_CP_6773_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/Update/ca
      -- 
    ca_7635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2912_inst_ack_1, ack => convTransposeD_CP_6773_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/$exit
      -- CP-element group 104: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/$exit
      -- CP-element group 104: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2912/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_req
      -- 
    phi_stmt_2907_req_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2907_req_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(104), ack => phi_stmt_2907_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(102) & convTransposeD_CP_6773_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/ra
      -- 
    ra_7653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2918_inst_ack_0, ack => convTransposeD_CP_6773_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/ca
      -- 
    ca_7658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2918_inst_ack_1, ack => convTransposeD_CP_6773_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/$exit
      -- CP-element group 107: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/$exit
      -- CP-element group 107: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_req
      -- 
    phi_stmt_2913_req_7659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2913_req_7659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(107), ack => phi_stmt_2913_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(105) & convTransposeD_CP_6773_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2580/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(101) & convTransposeD_CP_6773_elements(104) & convTransposeD_CP_6773_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Sample/ra
      -- 
    ra_7679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2903_inst_ack_0, ack => convTransposeD_CP_6773_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/Update/ca
      -- 
    ca_7684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2903_inst_ack_1, ack => convTransposeD_CP_6773_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/$exit
      -- CP-element group 111: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/$exit
      -- CP-element group 111: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_sources/type_cast_2903/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2900/phi_stmt_2900_req
      -- 
    phi_stmt_2900_req_7685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2900_req_7685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(111), ack => phi_stmt_2900_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(109) & convTransposeD_CP_6773_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Sample/ra
      -- 
    ra_7702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2910_inst_ack_0, ack => convTransposeD_CP_6773_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/Update/ca
      -- 
    ca_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2910_inst_ack_1, ack => convTransposeD_CP_6773_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/$exit
      -- CP-element group 114: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/$exit
      -- CP-element group 114: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_sources/type_cast_2910/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2907/phi_stmt_2907_req
      -- 
    phi_stmt_2907_req_7708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2907_req_7708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(114), ack => phi_stmt_2907_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(112) & convTransposeD_CP_6773_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/ra
      -- 
    ra_7725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2916_inst_ack_0, ack => convTransposeD_CP_6773_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/ca
      -- 
    ca_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2916_inst_ack_1, ack => convTransposeD_CP_6773_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/$exit
      -- CP-element group 117: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/$exit
      -- CP-element group 117: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_req
      -- 
    phi_stmt_2913_req_7731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2913_req_7731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(117), ack => phi_stmt_2913_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(115) & convTransposeD_CP_6773_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2580/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(111) & convTransposeD_CP_6773_elements(114) & convTransposeD_CP_6773_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2580/merge_stmt_2899_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2580/merge_stmt_2899_PhiAck/$entry
      -- 
    convTransposeD_CP_6773_elements(119) <= OrReduce(convTransposeD_CP_6773_elements(108) & convTransposeD_CP_6773_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2580/merge_stmt_2899_PhiAck/phi_stmt_2900_ack
      -- 
    phi_stmt_2900_ack_7736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2900_ack_0, ack => convTransposeD_CP_6773_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2580/merge_stmt_2899_PhiAck/phi_stmt_2907_ack
      -- 
    phi_stmt_2907_ack_7737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2907_ack_0, ack => convTransposeD_CP_6773_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2580/merge_stmt_2899_PhiAck/phi_stmt_2913_ack
      -- 
    phi_stmt_2913_ack_7738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2913_ack_0, ack => convTransposeD_CP_6773_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2580/merge_stmt_2899_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(120) & convTransposeD_CP_6773_elements(121) & convTransposeD_CP_6773_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2823_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2823_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2800_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2800_scaled : std_logic_vector(13 downto 0);
    signal add103_2858 : std_logic_vector(15 downto 0);
    signal add32_2659 : std_logic_vector(15 downto 0);
    signal add50_2665 : std_logic_vector(15 downto 0);
    signal add63_2676 : std_logic_vector(15 downto 0);
    signal add82_2776 : std_logic_vector(63 downto 0);
    signal add84_2786 : std_logic_vector(63 downto 0);
    signal add96_2840 : std_logic_vector(31 downto 0);
    signal add_2632 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2734 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2801_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2801_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2801_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2801_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2801_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2801_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2824_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2803 : std_logic_vector(31 downto 0);
    signal arrayidx92_2826 : std_logic_vector(31 downto 0);
    signal call11_2601 : std_logic_vector(15 downto 0);
    signal call13_2604 : std_logic_vector(15 downto 0);
    signal call14_2607 : std_logic_vector(15 downto 0);
    signal call15_2610 : std_logic_vector(15 downto 0);
    signal call16_2623 : std_logic_vector(15 downto 0);
    signal call18_2635 : std_logic_vector(15 downto 0);
    signal call1_2586 : std_logic_vector(15 downto 0);
    signal call20_2638 : std_logic_vector(15 downto 0);
    signal call22_2641 : std_logic_vector(15 downto 0);
    signal call3_2589 : std_logic_vector(15 downto 0);
    signal call5_2592 : std_logic_vector(15 downto 0);
    signal call7_2595 : std_logic_vector(15 downto 0);
    signal call9_2598 : std_logic_vector(15 downto 0);
    signal call_2583 : std_logic_vector(15 downto 0);
    signal cmp111_2871 : std_logic_vector(0 downto 0);
    signal cmp121_2892 : std_logic_vector(0 downto 0);
    signal cmp_2845 : std_logic_vector(0 downto 0);
    signal conv17_2627 : std_logic_vector(31 downto 0);
    signal conv70_2758 : std_logic_vector(63 downto 0);
    signal conv73_2685 : std_logic_vector(63 downto 0);
    signal conv75_2762 : std_logic_vector(63 downto 0);
    signal conv78_2689 : std_logic_vector(63 downto 0);
    signal conv80_2766 : std_logic_vector(63 downto 0);
    signal conv95_2834 : std_logic_vector(31 downto 0);
    signal conv99_2693 : std_logic_vector(31 downto 0);
    signal conv_2614 : std_logic_vector(31 downto 0);
    signal idxprom91_2819 : std_logic_vector(63 downto 0);
    signal idxprom_2796 : std_logic_vector(63 downto 0);
    signal inc115_2875 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2880 : std_logic_vector(15 downto 0);
    signal inc_2866 : std_logic_vector(15 downto 0);
    signal indvar_2696 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2925 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2913 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2717 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2907 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2710 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2887 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2900 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2703 : std_logic_vector(15 downto 0);
    signal mul59_2749 : std_logic_vector(15 downto 0);
    signal mul81_2771 : std_logic_vector(63 downto 0);
    signal mul83_2781 : std_logic_vector(63 downto 0);
    signal mul_2739 : std_logic_vector(15 downto 0);
    signal ptr_deref_2806_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2806_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2806_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2806_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2806_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2828_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2828_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2828_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2828_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2828_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2828_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2620 : std_logic_vector(31 downto 0);
    signal shr135_2648 : std_logic_vector(15 downto 0);
    signal shr31136_2654 : std_logic_vector(15 downto 0);
    signal shr86_2792 : std_logic_vector(31 downto 0);
    signal shr90_2813 : std_logic_vector(63 downto 0);
    signal sub53_2744 : std_logic_vector(15 downto 0);
    signal sub66_2681 : std_logic_vector(15 downto 0);
    signal sub67_2754 : std_logic_vector(15 downto 0);
    signal sub_2670 : std_logic_vector(15 downto 0);
    signal tmp1_2729 : std_logic_vector(31 downto 0);
    signal tmp88_2807 : std_logic_vector(63 downto 0);
    signal type_cast_2618_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2646_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2663_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2674_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2700_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2702_wire : std_logic_vector(31 downto 0);
    signal type_cast_2707_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2709_wire : std_logic_vector(15 downto 0);
    signal type_cast_2714_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2716_wire : std_logic_vector(15 downto 0);
    signal type_cast_2720_wire : std_logic_vector(15 downto 0);
    signal type_cast_2722_wire : std_logic_vector(15 downto 0);
    signal type_cast_2727_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2790_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2811_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2856_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2864_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2884_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2903_wire : std_logic_vector(15 downto 0);
    signal type_cast_2906_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2910_wire : std_logic_vector(15 downto 0);
    signal type_cast_2912_wire : std_logic_vector(15 downto 0);
    signal type_cast_2916_wire : std_logic_vector(15 downto 0);
    signal type_cast_2918_wire : std_logic_vector(15 downto 0);
    signal type_cast_2923_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2931_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2801_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2801_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2801_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2801_resized_base_address <= "00000000000000";
    array_obj_ref_2824_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2824_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2824_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2824_resized_base_address <= "00000000000000";
    ptr_deref_2806_word_offset_0 <= "00000000000000";
    ptr_deref_2828_word_offset_0 <= "00000000000000";
    type_cast_2618_wire_constant <= "00000000000000000000000000010000";
    type_cast_2646_wire_constant <= "0000000000000010";
    type_cast_2652_wire_constant <= "0000000000000001";
    type_cast_2663_wire_constant <= "1111111111111111";
    type_cast_2674_wire_constant <= "1111111111111111";
    type_cast_2700_wire_constant <= "00000000000000000000000000000000";
    type_cast_2707_wire_constant <= "0000000000000000";
    type_cast_2714_wire_constant <= "0000000000000000";
    type_cast_2727_wire_constant <= "00000000000000000000000000000100";
    type_cast_2790_wire_constant <= "00000000000000000000000000000010";
    type_cast_2811_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2817_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2838_wire_constant <= "00000000000000000000000000000100";
    type_cast_2856_wire_constant <= "0000000000000100";
    type_cast_2864_wire_constant <= "0000000000000001";
    type_cast_2884_wire_constant <= "0000000000000000";
    type_cast_2906_wire_constant <= "0000000000000000";
    type_cast_2923_wire_constant <= "00000000000000000000000000000001";
    type_cast_2931_wire_constant <= "0000000000000001";
    phi_stmt_2696: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2700_wire_constant & type_cast_2702_wire;
      req <= phi_stmt_2696_req_0 & phi_stmt_2696_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2696",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2696_ack_0,
          idata => idata,
          odata => indvar_2696,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2696
    phi_stmt_2703: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2707_wire_constant & type_cast_2709_wire;
      req <= phi_stmt_2703_req_0 & phi_stmt_2703_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2703",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2703_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2703,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2703
    phi_stmt_2710: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2714_wire_constant & type_cast_2716_wire;
      req <= phi_stmt_2710_req_0 & phi_stmt_2710_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2710",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2710_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2710,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2710
    phi_stmt_2717: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2720_wire & type_cast_2722_wire;
      req <= phi_stmt_2717_req_0 & phi_stmt_2717_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2717",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2717_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2717,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2717
    phi_stmt_2900: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2903_wire & type_cast_2906_wire_constant;
      req <= phi_stmt_2900_req_0 & phi_stmt_2900_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2900",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2900_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2900,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2900
    phi_stmt_2907: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2910_wire & type_cast_2912_wire;
      req <= phi_stmt_2907_req_0 & phi_stmt_2907_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2907",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2907_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2907,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2907
    phi_stmt_2913: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2916_wire & type_cast_2918_wire;
      req <= phi_stmt_2913_req_0 & phi_stmt_2913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2913",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2913_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2913
    -- flow-through select operator MUX_2886_inst
    input_dim1x_x2_2887 <= type_cast_2884_wire_constant when (cmp111_2871(0) /=  '0') else inc_2866;
    addr_of_2802_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2802_final_reg_req_0;
      addr_of_2802_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2802_final_reg_req_1;
      addr_of_2802_final_reg_ack_1<= rack(0);
      addr_of_2802_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2802_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2801_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2825_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2825_final_reg_req_0;
      addr_of_2825_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2825_final_reg_req_1;
      addr_of_2825_final_reg_ack_1<= rack(0);
      addr_of_2825_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2825_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2824_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2613_inst_req_0;
      type_cast_2613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2613_inst_req_1;
      type_cast_2613_inst_ack_1<= rack(0);
      type_cast_2613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2626_inst_req_0;
      type_cast_2626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2626_inst_req_1;
      type_cast_2626_inst_ack_1<= rack(0);
      type_cast_2626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2684_inst_req_0;
      type_cast_2684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2684_inst_req_1;
      type_cast_2684_inst_ack_1<= rack(0);
      type_cast_2684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2688_inst_req_0;
      type_cast_2688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2688_inst_req_1;
      type_cast_2688_inst_ack_1<= rack(0);
      type_cast_2688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2638,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2692_inst_req_0;
      type_cast_2692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2692_inst_req_1;
      type_cast_2692_inst_ack_1<= rack(0);
      type_cast_2692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2702_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2702_inst_req_0;
      type_cast_2702_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2702_inst_req_1;
      type_cast_2702_inst_ack_1<= rack(0);
      type_cast_2702_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2702_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2925,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2702_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2709_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2716_inst_req_0;
      type_cast_2716_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2716_inst_req_1;
      type_cast_2716_inst_ack_1<= rack(0);
      type_cast_2716_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2907,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2716_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2720_inst_req_0;
      type_cast_2720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2720_inst_req_1;
      type_cast_2720_inst_ack_1<= rack(0);
      type_cast_2720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2720_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2722_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2757_inst_req_0;
      type_cast_2757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2757_inst_req_1;
      type_cast_2757_inst_ack_1<= rack(0);
      type_cast_2757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2761_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2761_inst_req_0;
      type_cast_2761_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2761_inst_req_1;
      type_cast_2761_inst_ack_1<= rack(0);
      type_cast_2761_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2761_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2762,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2765_inst_req_0;
      type_cast_2765_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2765_inst_req_1;
      type_cast_2765_inst_ack_1<= rack(0);
      type_cast_2765_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2744,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2795_inst_req_0;
      type_cast_2795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2795_inst_req_1;
      type_cast_2795_inst_ack_1<= rack(0);
      type_cast_2795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2833_inst_req_0;
      type_cast_2833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2833_inst_req_1;
      type_cast_2833_inst_ack_1<= rack(0);
      type_cast_2833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2874_inst_req_0;
      type_cast_2874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2874_inst_req_1;
      type_cast_2874_inst_ack_1<= rack(0);
      type_cast_2874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2871,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2903_inst_req_0;
      type_cast_2903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2903_inst_req_1;
      type_cast_2903_inst_ack_1<= rack(0);
      type_cast_2903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2858,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2903_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2910_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2910_inst_req_0;
      type_cast_2910_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2910_inst_req_1;
      type_cast_2910_inst_ack_1<= rack(0);
      type_cast_2910_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2910_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2910_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2912_inst_req_0;
      type_cast_2912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2912_inst_req_1;
      type_cast_2912_inst_ack_1<= rack(0);
      type_cast_2912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2887,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2912_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2916_inst_req_0;
      type_cast_2916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2916_inst_req_1;
      type_cast_2916_inst_ack_1<= rack(0);
      type_cast_2916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2717,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2916_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2918_inst_req_0;
      type_cast_2918_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2918_inst_req_1;
      type_cast_2918_inst_ack_1<= rack(0);
      type_cast_2918_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2918_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2918_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2801_index_1_rename
    process(R_idxprom_2800_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2800_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2800_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2801_index_1_resize
    process(idxprom_2796) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2796;
      ov := iv(13 downto 0);
      R_idxprom_2800_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2801_root_address_inst
    process(array_obj_ref_2801_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2801_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2801_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2824_index_1_rename
    process(R_idxprom91_2823_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2823_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2823_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2824_index_1_resize
    process(idxprom91_2819) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2819;
      ov := iv(13 downto 0);
      R_idxprom91_2823_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2824_root_address_inst
    process(array_obj_ref_2824_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2824_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2824_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2806_addr_0
    process(ptr_deref_2806_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2806_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2806_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2806_base_resize
    process(arrayidx87_2803) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2803;
      ov := iv(13 downto 0);
      ptr_deref_2806_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2806_gather_scatter
    process(ptr_deref_2806_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2806_data_0;
      ov(63 downto 0) := iv;
      tmp88_2807 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2806_root_address_inst
    process(ptr_deref_2806_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2806_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2806_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2828_addr_0
    process(ptr_deref_2828_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2828_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2828_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2828_base_resize
    process(arrayidx92_2826) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2826;
      ov := iv(13 downto 0);
      ptr_deref_2828_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2828_gather_scatter
    process(tmp88_2807) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2807;
      ov(63 downto 0) := iv;
      ptr_deref_2828_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2828_root_address_inst
    process(ptr_deref_2828_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2828_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2828_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2846_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2845;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2846_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2846_branch_req_0,
          ack0 => if_stmt_2846_branch_ack_0,
          ack1 => if_stmt_2846_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2893_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2892;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2893_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2893_branch_req_0,
          ack0 => if_stmt_2893_branch_ack_0,
          ack1 => if_stmt_2893_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2658_inst
    process(shr135_2648, shr31136_2654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2648, shr31136_2654, tmp_var);
      add32_2659 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2664_inst
    process(call7_2595) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2595, type_cast_2663_wire_constant, tmp_var);
      add50_2665 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2675_inst
    process(call9_2598) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2598, type_cast_2674_wire_constant, tmp_var);
      add63_2676 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2743_inst
    process(sub_2670, mul_2739) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2670, mul_2739, tmp_var);
      sub53_2744 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2753_inst
    process(sub66_2681, mul59_2749) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2681, mul59_2749, tmp_var);
      sub67_2754 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2857_inst
    process(input_dim2x_x1_2703) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2703, type_cast_2856_wire_constant, tmp_var);
      add103_2858 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2865_inst
    process(input_dim1x_x1_2710) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2710, type_cast_2864_wire_constant, tmp_var);
      inc_2866 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2879_inst
    process(inc115_2875, input_dim0x_x2_2717) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2875, input_dim0x_x2_2717, tmp_var);
      inc115x_xinput_dim0x_x2_2880 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2733_inst
    process(add_2632, tmp1_2729) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2632, tmp1_2729, tmp_var);
      add_src_0x_x0_2734 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2839_inst
    process(conv95_2834) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2834, type_cast_2838_wire_constant, tmp_var);
      add96_2840 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2924_inst
    process(indvar_2696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2696, type_cast_2923_wire_constant, tmp_var);
      indvarx_xnext_2925 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2775_inst
    process(mul81_2771, conv75_2762) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2771, conv75_2762, tmp_var);
      add82_2776 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2785_inst
    process(mul83_2781, conv70_2758) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2781, conv70_2758, tmp_var);
      add84_2786 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2818_inst
    process(shr90_2813) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2813, type_cast_2817_wire_constant, tmp_var);
      idxprom91_2819 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2870_inst
    process(inc_2866, call1_2586) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2866, call1_2586, tmp_var);
      cmp111_2871 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2891_inst
    process(inc115x_xinput_dim0x_x2_2880, call_2583) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2880, call_2583, tmp_var);
      cmp121_2892 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2647_inst
    process(call_2583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2583, type_cast_2646_wire_constant, tmp_var);
      shr135_2648 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2653_inst
    process(call_2583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2583, type_cast_2652_wire_constant, tmp_var);
      shr31136_2654 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2791_inst
    process(add_src_0x_x0_2734) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2734, type_cast_2790_wire_constant, tmp_var);
      shr86_2792 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2812_inst
    process(add84_2786) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2786, type_cast_2811_wire_constant, tmp_var);
      shr90_2813 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2738_inst
    process(input_dim0x_x2_2717, call13_2604) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2717, call13_2604, tmp_var);
      mul_2739 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2748_inst
    process(input_dim1x_x1_2710, call13_2604) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2710, call13_2604, tmp_var);
      mul59_2749 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2728_inst
    process(indvar_2696) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2696, type_cast_2727_wire_constant, tmp_var);
      tmp1_2729 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2770_inst
    process(conv80_2766, conv78_2689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2766, conv78_2689, tmp_var);
      mul81_2771 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2780_inst
    process(add82_2776, conv73_2685) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2776, conv73_2685, tmp_var);
      mul83_2781 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2631_inst
    process(shl_2620, conv17_2627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2620, conv17_2627, tmp_var);
      add_2632 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2619_inst
    process(conv_2614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2614, type_cast_2618_wire_constant, tmp_var);
      shl_2620 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2669_inst
    process(add50_2665, call14_2607) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2665, call14_2607, tmp_var);
      sub_2670 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2680_inst
    process(add63_2676, call14_2607) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2676, call14_2607, tmp_var);
      sub66_2681 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2844_inst
    process(add96_2840, conv99_2693) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2840, conv99_2693, tmp_var);
      cmp_2845 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2801_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2800_scaled;
      array_obj_ref_2801_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2801_index_offset_req_0;
      array_obj_ref_2801_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2801_index_offset_req_1;
      array_obj_ref_2801_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2824_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2823_scaled;
      array_obj_ref_2824_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2824_index_offset_req_0;
      array_obj_ref_2824_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2824_index_offset_req_1;
      array_obj_ref_2824_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2806_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2806_load_0_req_0;
      ptr_deref_2806_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2806_load_0_req_1;
      ptr_deref_2806_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2806_word_address_0;
      ptr_deref_2806_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2828_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2828_store_0_req_0;
      ptr_deref_2828_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2828_store_0_req_1;
      ptr_deref_2828_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2828_word_address_0;
      data_in <= ptr_deref_2828_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2582_inst RPIPE_Block3_start_2585_inst RPIPE_Block3_start_2588_inst RPIPE_Block3_start_2591_inst RPIPE_Block3_start_2594_inst RPIPE_Block3_start_2597_inst RPIPE_Block3_start_2600_inst RPIPE_Block3_start_2603_inst RPIPE_Block3_start_2606_inst RPIPE_Block3_start_2609_inst RPIPE_Block3_start_2622_inst RPIPE_Block3_start_2634_inst RPIPE_Block3_start_2637_inst RPIPE_Block3_start_2640_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2582_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2585_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2588_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2591_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2594_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2597_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2600_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2603_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2606_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2609_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2622_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2634_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2637_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2640_inst_req_0;
      RPIPE_Block3_start_2582_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2585_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2588_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2591_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2594_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2597_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2600_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2603_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2606_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2609_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2622_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2634_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2637_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2640_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2582_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2585_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2588_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2591_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2594_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2597_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2600_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2603_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2606_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2609_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2622_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2634_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2637_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2640_inst_req_1;
      RPIPE_Block3_start_2582_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2585_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2588_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2591_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2594_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2597_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2600_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2603_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2606_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2609_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2622_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2634_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2637_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2640_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2583 <= data_out(223 downto 208);
      call1_2586 <= data_out(207 downto 192);
      call3_2589 <= data_out(191 downto 176);
      call5_2592 <= data_out(175 downto 160);
      call7_2595 <= data_out(159 downto 144);
      call9_2598 <= data_out(143 downto 128);
      call11_2601 <= data_out(127 downto 112);
      call13_2604 <= data_out(111 downto 96);
      call14_2607 <= data_out(95 downto 80);
      call15_2610 <= data_out(79 downto 64);
      call16_2623 <= data_out(63 downto 48);
      call18_2635 <= data_out(47 downto 32);
      call20_2638 <= data_out(31 downto 16);
      call22_2641 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2929_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2929_inst_req_0;
      WPIPE_Block3_done_2929_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2929_inst_req_1;
      WPIPE_Block3_done_2929_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2931_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_28_load_0_req_1 : boolean;
  signal LOAD_count_28_load_0_ack_1 : boolean;
  signal LOAD_count_28_load_0_req_0 : boolean;
  signal LOAD_count_28_load_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_update_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/rr
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_sample_completed_
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/ra
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_ack
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_29/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_update_completed_
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_28_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_28_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_28_word_address_0 <= "0";
    -- equivalence LOAD_count_28_gather_scatter
    process(LOAD_count_28_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_28_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_28_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_28_load_0_req_0;
      LOAD_count_28_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_28_load_0_req_1;
      LOAD_count_28_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_28_word_address_0;
      LOAD_count_28_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
