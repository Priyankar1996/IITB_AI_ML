-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_45_branch_req_0 : boolean;
  signal phi_stmt_47_req_0 : boolean;
  signal phi_stmt_47_req_1 : boolean;
  signal phi_stmt_47_ack_0 : boolean;
  signal n_address_281_49_buf_req_0 : boolean;
  signal n_address_281_49_buf_ack_0 : boolean;
  signal n_address_281_49_buf_req_1 : boolean;
  signal n_address_281_49_buf_ack_1 : boolean;
  signal phi_stmt_52_req_1 : boolean;
  signal phi_stmt_52_req_0 : boolean;
  signal phi_stmt_52_ack_0 : boolean;
  signal n_word_start_270_57_buf_req_0 : boolean;
  signal n_word_start_270_57_buf_ack_0 : boolean;
  signal n_word_start_270_57_buf_req_1 : boolean;
  signal n_word_start_270_57_buf_ack_1 : boolean;
  signal n_winr_210_71_buf_req_0 : boolean;
  signal n_winr_210_71_buf_ack_0 : boolean;
  signal n_winr_210_71_buf_req_1 : boolean;
  signal phi_stmt_58_req_0 : boolean;
  signal phi_stmt_58_req_1 : boolean;
  signal phi_stmt_58_ack_0 : boolean;
  signal n_left_289_60_buf_req_0 : boolean;
  signal n_left_289_60_buf_ack_0 : boolean;
  signal n_left_289_60_buf_req_1 : boolean;
  signal n_left_289_60_buf_ack_1 : boolean;
  signal nl_start_36_61_buf_req_0 : boolean;
  signal nl_start_36_61_buf_ack_0 : boolean;
  signal nl_start_36_61_buf_req_1 : boolean;
  signal nl_start_36_61_buf_ack_1 : boolean;
  signal phi_stmt_62_req_0 : boolean;
  signal phi_stmt_62_req_1 : boolean;
  signal phi_stmt_62_ack_0 : boolean;
  signal n_blk_309_64_buf_req_0 : boolean;
  signal n_blk_309_64_buf_ack_0 : boolean;
  signal n_blk_309_64_buf_req_1 : boolean;
  signal n_blk_309_64_buf_ack_1 : boolean;
  signal type_cast_66_inst_req_0 : boolean;
  signal type_cast_66_inst_ack_0 : boolean;
  signal type_cast_66_inst_req_1 : boolean;
  signal type_cast_66_inst_ack_1 : boolean;
  signal phi_stmt_67_req_1 : boolean;
  signal phi_stmt_67_req_0 : boolean;
  signal phi_stmt_67_ack_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_req_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_ack_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_req_1 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_ack_1 : boolean;
  signal n_winr_210_71_buf_ack_1 : boolean;
  signal phi_stmt_72_req_0 : boolean;
  signal phi_stmt_72_req_1 : boolean;
  signal phi_stmt_72_ack_0 : boolean;
  signal n_col_223_74_buf_req_0 : boolean;
  signal n_col_223_74_buf_ack_0 : boolean;
  signal n_col_223_74_buf_req_1 : boolean;
  signal n_col_223_74_buf_ack_1 : boolean;
  signal phi_stmt_77_req_0 : boolean;
  signal phi_stmt_77_req_1 : boolean;
  signal phi_stmt_77_ack_0 : boolean;
  signal n_row_235_79_buf_req_0 : boolean;
  signal n_row_235_79_buf_ack_0 : boolean;
  signal n_row_235_79_buf_req_1 : boolean;
  signal n_row_235_79_buf_ack_1 : boolean;
  signal array_obj_ref_134_index_offset_req_0 : boolean;
  signal array_obj_ref_134_index_offset_ack_0 : boolean;
  signal array_obj_ref_134_index_offset_req_1 : boolean;
  signal array_obj_ref_134_index_offset_ack_1 : boolean;
  signal addr_of_135_final_reg_req_0 : boolean;
  signal addr_of_135_final_reg_ack_0 : boolean;
  signal addr_of_135_final_reg_req_1 : boolean;
  signal addr_of_135_final_reg_ack_1 : boolean;
  signal ptr_deref_139_load_0_req_0 : boolean;
  signal ptr_deref_139_load_0_ack_0 : boolean;
  signal ptr_deref_139_load_0_req_1 : boolean;
  signal ptr_deref_139_load_0_ack_1 : boolean;
  signal slice_143_inst_req_0 : boolean;
  signal slice_143_inst_ack_0 : boolean;
  signal slice_143_inst_req_1 : boolean;
  signal slice_143_inst_ack_1 : boolean;
  signal slice_147_inst_req_0 : boolean;
  signal slice_147_inst_ack_0 : boolean;
  signal slice_147_inst_req_1 : boolean;
  signal slice_147_inst_ack_1 : boolean;
  signal slice_151_inst_req_0 : boolean;
  signal slice_151_inst_ack_0 : boolean;
  signal slice_151_inst_req_1 : boolean;
  signal slice_151_inst_ack_1 : boolean;
  signal slice_155_inst_req_0 : boolean;
  signal slice_155_inst_ack_0 : boolean;
  signal slice_155_inst_req_1 : boolean;
  signal slice_155_inst_ack_1 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_req_0 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_ack_0 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_req_1 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_161_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_161_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_161_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_161_inst_ack_1 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_req_0 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_ack_0 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_req_1 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_168_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_168_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_168_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_168_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_175_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_175_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_175_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_175_inst_ack_1 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_req_0 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_ack_0 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_req_1 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_182_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_182_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_182_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_182_inst_ack_1 : boolean;
  signal do_while_stmt_45_branch_ack_0 : boolean;
  signal do_while_stmt_45_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_27/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/branch_block_stmt_27__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44__exit__
      -- CP-element group 0: 	 branch_block_stmt_27/do_while_stmt_45__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_27/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/branch_block_stmt_27__exit__
      -- CP-element group 1: 	 branch_block_stmt_27/do_while_stmt_45__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_27/do_while_stmt_45/$entry
      -- CP-element group 2: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_27/do_while_stmt_45/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/condition_done
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_27/do_while_stmt_45/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	117 
    -- CP-element group 7: 	99 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	78 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	59 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	119 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	80 
    -- CP-element group 8: 	101 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	61 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	113 
    -- CP-element group 9: 	112 
    -- CP-element group 9: 	94 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	130 
    -- CP-element group 9: 	131 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	73 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	203 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_45_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(14) & access_T_CP_0_elements(203);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	130 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	114 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	55 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(112) & access_T_CP_0_elements(93) & access_T_CP_0_elements(130) & access_T_CP_0_elements(15) & access_T_CP_0_elements(34) & access_T_CP_0_elements(53) & access_T_CP_0_elements(72) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	115 
    -- CP-element group 12: 	96 
    -- CP-element group 12: 	132 
    -- CP-element group 12: 	75 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	56 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	112 
    -- CP-element group 12: 	93 
    -- CP-element group 12: 	130 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	72 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(115) & access_T_CP_0_elements(96) & access_T_CP_0_elements(132) & access_T_CP_0_elements(75) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	113 
    -- CP-element group 13: 	94 
    -- CP-element group 13: 	131 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	73 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	76 
    -- CP-element group 13: 	97 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	57 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(113) & access_T_CP_0_elements(94) & access_T_CP_0_elements(131) & access_T_CP_0_elements(16) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54) & access_T_CP_0_elements(73);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	77 
    -- CP-element group 14: 	98 
    -- CP-element group 14: 	116 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(98) & access_T_CP_0_elements(116) & access_T_CP_0_elements(134) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: 	151 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_134_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_sample_req_ps
      -- 
    phi_stmt_47_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_47_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_47_req_0); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_sample_req_ps
      -- 
    phi_stmt_47_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_47_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_47_req_1); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_phi_mux_ack_ps
      -- 
    phi_stmt_47_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_47_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Sample/req
      -- 
    req_63_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_63_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(26), ack => n_address_281_49_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_update_start_
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Update/req
      -- 
    req_68_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_68_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(27), ack => n_address_281_49_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Sample/ack
      -- 
    ack_64_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_281_49_buf_ack_0, ack => access_T_CP_0_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_49_Update/ack
      -- 
    ack_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_281_49_buf_ack_1, ack => access_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_update_start_
      -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_update_completed__ps
      -- 
    access_T_CP_0_elements(32) <= access_T_CP_0_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_51_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(31), ack => access_T_CP_0_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	177 
    -- CP-element group 35: 	184 
    -- CP-element group 35: 	191 
    -- CP-element group 35: 	198 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	175 
    -- CP-element group 39: 	182 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	189 
    -- CP-element group 39: 	196 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_sample_req_ps
      -- 
    phi_stmt_52_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_52_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_52_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_sample_req_ps
      -- 
    phi_stmt_52_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_52_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_52_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_phi_mux_ack_ps
      -- 
    phi_stmt_52_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_52_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(49), ack => n_word_start_270_57_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_start_
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(50), ack => n_word_start_270_57_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_270_57_buf_ack_0, ack => access_T_CP_0_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_270_57_buf_ack_1, ack => access_T_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_start_
      -- 
    access_T_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_start_
      -- 
    access_T_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_sample_req_ps
      -- 
    phi_stmt_58_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_58_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_58_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_sample_req_ps
      -- 
    phi_stmt_58_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_58_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_58_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_phi_mux_ack_ps
      -- 
    phi_stmt_58_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_58_ack_0, ack => access_T_CP_0_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => n_left_289_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_start_
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(65), ack => n_left_289_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_289_60_buf_ack_0, ack => access_T_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_289_60_buf_ack_1, ack => access_T_CP_0_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => nl_start_36_61_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_start_
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => nl_start_36_61_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_36_61_buf_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_36_61_buf_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	12 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	11 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_start_
      -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	184 
    -- CP-element group 73: 	191 
    -- CP-element group 73: 	198 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	13 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_start_
      -- 
    access_T_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	11 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(11);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	12 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	13 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_start__ps
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(13);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	182 
    -- CP-element group 77: 	14 
    -- CP-element group 77: 	189 
    -- CP-element group 77: 	196 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	7 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(7);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_sample_req
      -- CP-element group 79: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_sample_req_ps
      -- 
    phi_stmt_62_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_62_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_62_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	8 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_trigger
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(8);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_sample_req
      -- CP-element group 81: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_sample_req_ps
      -- 
    phi_stmt_62_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_62_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => phi_stmt_62_req_1); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_phi_mux_ack
      -- CP-element group 82: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_phi_mux_ack_ps
      -- 
    phi_stmt_62_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_62_ack_0, ack => access_T_CP_0_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_start__ps
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/req
      -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => n_blk_309_64_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_start__ps
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_start_
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/req
      -- 
    req_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => n_blk_309_64_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/ack
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_309_64_buf_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/ack
      -- 
    ack_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_309_64_buf_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/rr
      -- 
    rr_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => type_cast_66_inst_req_0); -- 
    access_T_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(87) & access_T_CP_0_elements(91);
      gj_access_T_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_start_
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/cr
      -- 
    cr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(90), ack => type_cast_66_inst_req_1); -- 
    access_T_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(88) & access_T_CP_0_elements(92);
      gj_access_T_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/ra
      -- 
    ra_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_0, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/ca
      -- 
    ca_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_1, ack => access_T_CP_0_elements(92)); -- 
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	11 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_start_
      -- 
    access_T_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	9 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	13 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_start_
      -- 
    access_T_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(98);
      gj_access_T_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(11);
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	12 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	13 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_start__ps
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(13);
    -- CP-element group 98:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	14 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	94 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	7 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(7);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_sample_req
      -- CP-element group 100: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_sample_req_ps
      -- 
    phi_stmt_67_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_67_req_1); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	8 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_trigger
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(8);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_sample_req
      -- CP-element group 102: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_sample_req_ps
      -- 
    phi_stmt_67_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => phi_stmt_67_req_0); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_phi_mux_ack
      -- CP-element group 103: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_phi_mux_ack_ps
      -- 
    phi_stmt_67_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_67_ack_0, ack => access_T_CP_0_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_start_
      -- 
    -- Element group access_T_CP_0_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_completed__ps
      -- 
    access_T_CP_0_elements(106) <= access_T_CP_0_elements(107);
    -- CP-element group 107:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	106 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(107) is a control-delay.
    cp_element_107_delay: control_delay_element  generic map(name => " 107_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(105), ack => access_T_CP_0_elements(107), clk => clk, reset =>reset);
    -- CP-element group 108:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/req
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_start__ps
      -- 
    req_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(108), ack => n_winr_210_71_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_start_
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/req
      -- 
    req_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(109), ack => n_winr_210_71_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_completed__ps
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/ack
      -- 
    ack_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_210_71_buf_ack_0, ack => access_T_CP_0_elements(110)); -- 
    -- CP-element group 111:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_completed__ps
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/ack
      -- 
    ack_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_210_71_buf_ack_1, ack => access_T_CP_0_elements(111)); -- 
    -- CP-element group 112:  join  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	9 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	12 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	11 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_start_
      -- 
    access_T_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	9 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	116 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	13 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_start_
      -- 
    access_T_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(116);
      gj_access_T_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	11 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(11);
    -- CP-element group 115:  join  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	12 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	14 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	113 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(116) is bound as output of CP function.
    -- CP-element group 117:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	7 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_trigger
      -- 
    access_T_CP_0_elements(117) <= access_T_CP_0_elements(7);
    -- CP-element group 118:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_sample_req
      -- CP-element group 118: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_sample_req_ps
      -- 
    phi_stmt_72_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(118), ack => phi_stmt_72_req_0); -- 
    -- Element group access_T_CP_0_elements(118) is bound as output of CP function.
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	8 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_trigger
      -- 
    access_T_CP_0_elements(119) <= access_T_CP_0_elements(8);
    -- CP-element group 120:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_sample_req
      -- CP-element group 120: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_sample_req_ps
      -- 
    phi_stmt_72_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(120), ack => phi_stmt_72_req_1); -- 
    -- Element group access_T_CP_0_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_phi_mux_ack
      -- CP-element group 121: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_phi_mux_ack_ps
      -- 
    phi_stmt_72_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_72_ack_0, ack => access_T_CP_0_elements(121)); -- 
    -- CP-element group 122:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_start__ps
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/req
      -- 
    req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(122), ack => n_col_223_74_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_start__ps
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_start_
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(123), ack => n_col_223_74_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_completed__ps
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/ack
      -- 
    ack_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_223_74_buf_ack_0, ack => access_T_CP_0_elements(124)); -- 
    -- CP-element group 125:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/ack
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_223_74_buf_ack_1, ack => access_T_CP_0_elements(125)); -- 
    -- CP-element group 126:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_start__ps
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_start__ps
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_start_
      -- 
    -- Element group access_T_CP_0_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_completed__ps
      -- 
    access_T_CP_0_elements(128) <= access_T_CP_0_elements(129);
    -- CP-element group 129:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	128 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(129) is a control-delay.
    cp_element_129_delay: control_delay_element  generic map(name => " 129_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(127), ack => access_T_CP_0_elements(129), clk => clk, reset =>reset);
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	12 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	11 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	9 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	134 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	13 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_start_
      -- 
    access_T_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	131 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_sample_req_ps
      -- 
    phi_stmt_77_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_77_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_77_req_0); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_sample_req_ps
      -- 
    phi_stmt_77_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_77_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_77_req_1); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_phi_mux_ack_ps
      -- 
    phi_stmt_77_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_77_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Sample/req
      -- 
    req_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(140), ack => n_row_235_79_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_update_start_
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Update/req
      -- 
    req_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(141), ack => n_row_235_79_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_sample_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Sample/ack
      -- 
    ack_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_235_79_buf_ack_0, ack => access_T_CP_0_elements(142)); -- 
    -- CP-element group 143:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_update_completed__ps
      -- CP-element group 143: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_79_Update/ack
      -- 
    ack_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_235_79_buf_ack_1, ack => access_T_CP_0_elements(143)); -- 
    -- CP-element group 144:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_update_start_
      -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_update_completed__ps
      -- 
    access_T_CP_0_elements(146) <= access_T_CP_0_elements(147);
    -- CP-element group 147:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_81_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(147) is a control-delay.
    cp_element_147_delay: control_delay_element  generic map(name => " 147_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(145), ack => access_T_CP_0_elements(147), clk => clk, reset =>reset);
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_135_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_update_start_
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_135_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_134_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	20 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_134_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_134_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_135_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_135_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_139_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	169 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_update_start_
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_139_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(173) & access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	171 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_143_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_update_start_
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_143_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_143_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_143_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_147_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_update_start_
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_147_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	156 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_151_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_update_start_
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_151_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	156 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_155_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_update_start_
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_155_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	156 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	39 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_157_delayed_14_0_157_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_update_start_
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_157_delayed_14_0_157_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	35 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_157_delayed_14_0_157_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_157_delayed_14_0_157_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	162 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_161_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(162) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	160 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_update_start_
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_161_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_161_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_161_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	77 
    -- CP-element group 182: 	39 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_161_delayed_14_0_164_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_update_start_
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_161_delayed_14_0_164_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	35 
    -- CP-element group 184: 	73 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_161_delayed_14_0_164_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_161_delayed_14_0_164_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	166 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_168_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(181) & access_T_CP_0_elements(185) & access_T_CP_0_elements(166) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_update_start_
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/req
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_168_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_168_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/ack
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_168_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	77 
    -- CP-element group 189: 	39 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_165_delayed_14_0_171_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_update_start_
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_165_delayed_14_0_171_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	35 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	73 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_165_delayed_14_0_171_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_165_delayed_14_0_171_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	170 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_175_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(170) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_update_start_
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_175_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_175_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_175_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	77 
    -- CP-element group 196: 	39 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_169_delayed_14_0_178_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(39) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_update_start_
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_169_delayed_14_0_178_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	35 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	73 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_169_delayed_14_0_178_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_169_delayed_14_0_178_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_182_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(174) & access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	172 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_update_start_
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_182_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_182_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_182_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(12) & access_T_CP_0_elements(151) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_45_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_45_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_27/do_while_stmt_45/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_45_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_45_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_47_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(29);
      access_T_CP_0_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(30);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(24) <= phi_mux_reqs(1);
      phi_stmt_47_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_47_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_52_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(51);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(52);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_52_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_52_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_58_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(67);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_58_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_58_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(55), 
          phi_sample_ack => access_T_CP_0_elements(56), 
          phi_update_req => access_T_CP_0_elements(57), 
          phi_update_ack => access_T_CP_0_elements(58), 
          phi_mux_ack => access_T_CP_0_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_62_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(80);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(92);
      access_T_CP_0_elements(81) <= phi_mux_reqs(1);
      phi_stmt_62_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_62_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(74), 
          phi_sample_ack => access_T_CP_0_elements(75), 
          phi_update_req => access_T_CP_0_elements(76), 
          phi_update_ack => access_T_CP_0_elements(77), 
          phi_mux_ack => access_T_CP_0_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_67_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(101);
      access_T_CP_0_elements(104)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(105)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(102) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(108)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(110);
      access_T_CP_0_elements(109)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(111);
      access_T_CP_0_elements(100) <= phi_mux_reqs(1);
      phi_stmt_67_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_67_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(95), 
          phi_sample_ack => access_T_CP_0_elements(96), 
          phi_update_req => access_T_CP_0_elements(97), 
          phi_update_ack => access_T_CP_0_elements(98), 
          phi_mux_ack => access_T_CP_0_elements(103), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_72_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(117);
      access_T_CP_0_elements(122)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(123)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(125);
      access_T_CP_0_elements(118) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(119);
      access_T_CP_0_elements(126)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(126);
      access_T_CP_0_elements(127)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(120) <= phi_mux_reqs(1);
      phi_stmt_72_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_72_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(114), 
          phi_sample_ack => access_T_CP_0_elements(115), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(116), 
          phi_mux_ack => access_T_CP_0_elements(121), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_77_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(136) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(138) <= phi_mux_reqs(1);
      phi_stmt_77_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_77_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_126_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_206_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_219_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_232_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_294_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_279_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_108_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_115_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_214_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_229_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_95_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_261_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_104_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_111_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_118_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_91_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_98_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_275_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_243_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_31_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_250_wire : std_logic_vector(31 downto 0);
    signal MUX_207_wire : std_logic_vector(15 downto 0);
    signal MUX_220_wire : std_logic_vector(15 downto 0);
    signal MUX_301_wire : std_logic_vector(15 downto 0);
    signal MUX_307_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_313_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_119_wire : std_logic_vector(0 downto 0);
    signal R_address_133_resized : std_logic_vector(13 downto 0);
    signal R_address_133_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_287_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_299_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_107_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_114_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_296_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_94_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_304_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_40_wire : std_logic_vector(0 downto 0);
    signal address_47 : std_logic_vector(63 downto 0);
    signal array_obj_ref_134_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_root_address : std_logic_vector(13 downto 0);
    signal c1_157_delayed_14_0_159 : std_logic_vector(0 downto 0);
    signal c1_87 : std_logic_vector(0 downto 0);
    signal c2_100 : std_logic_vector(0 downto 0);
    signal c2_161_delayed_14_0_166 : std_logic_vector(0 downto 0);
    signal c3_121 : std_logic_vector(0 downto 0);
    signal c3_165_delayed_14_0_173 : std_logic_vector(0 downto 0);
    signal c4_129 : std_logic_vector(0 downto 0);
    signal c4_169_delayed_14_0_180 : std_logic_vector(0 downto 0);
    signal col_72 : std_logic_vector(15 downto 0);
    signal col_done_199 : std_logic_vector(0 downto 0);
    signal fetch_addr_136 : std_logic_vector(31 downto 0);
    signal flag1_189 : std_logic_vector(0 downto 0);
    signal fn_blk_44 : std_logic_vector(15 downto 0);
    signal konst_103_wire_constant : std_logic_vector(1 downto 0);
    signal konst_106_wire_constant : std_logic_vector(15 downto 0);
    signal konst_110_wire_constant : std_logic_vector(1 downto 0);
    signal konst_113_wire_constant : std_logic_vector(15 downto 0);
    signal konst_117_wire_constant : std_logic_vector(1 downto 0);
    signal konst_127_wire_constant : std_logic_vector(15 downto 0);
    signal konst_203_wire_constant : std_logic_vector(15 downto 0);
    signal konst_205_wire_constant : std_logic_vector(15 downto 0);
    signal konst_216_wire_constant : std_logic_vector(15 downto 0);
    signal konst_218_wire_constant : std_logic_vector(15 downto 0);
    signal konst_231_wire_constant : std_logic_vector(15 downto 0);
    signal konst_260_wire_constant : std_logic_vector(31 downto 0);
    signal konst_268_wire_constant : std_logic_vector(1 downto 0);
    signal konst_274_wire_constant : std_logic_vector(31 downto 0);
    signal konst_278_wire_constant : std_logic_vector(63 downto 0);
    signal konst_295_wire_constant : std_logic_vector(15 downto 0);
    signal konst_297_wire_constant : std_logic_vector(15 downto 0);
    signal konst_303_wire_constant : std_logic_vector(15 downto 0);
    signal konst_306_wire_constant : std_logic_vector(15 downto 0);
    signal konst_39_wire_constant : std_logic_vector(15 downto 0);
    signal konst_42_wire_constant : std_logic_vector(15 downto 0);
    signal konst_85_wire_constant : std_logic_vector(1 downto 0);
    signal konst_90_wire_constant : std_logic_vector(1 downto 0);
    signal konst_93_wire_constant : std_logic_vector(15 downto 0);
    signal konst_97_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_33 : std_logic_vector(31 downto 0);
    signal n_address_281 : std_logic_vector(63 downto 0);
    signal n_address_281_49_buffered : std_logic_vector(63 downto 0);
    signal n_blk_309 : std_logic_vector(15 downto 0);
    signal n_blk_309_64_buffered : std_logic_vector(15 downto 0);
    signal n_col_223 : std_logic_vector(15 downto 0);
    signal n_col_223_74_buffered : std_logic_vector(15 downto 0);
    signal n_left_289 : std_logic_vector(15 downto 0);
    signal n_left_289_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_235 : std_logic_vector(15 downto 0);
    signal n_row_235_79_buffered : std_logic_vector(15 downto 0);
    signal n_winr_210 : std_logic_vector(15 downto 0);
    signal n_winr_210_71_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_270 : std_logic_vector(1 downto 0);
    signal n_word_start_270_57_buffered : std_logic_vector(1 downto 0);
    signal na1_245 : std_logic_vector(31 downto 0);
    signal na2_252 : std_logic_vector(31 downto 0);
    signal na3_257 : std_logic_vector(31 downto 0);
    signal na4_263 : std_logic_vector(15 downto 0);
    signal nl_start_36 : std_logic_vector(15 downto 0);
    signal nl_start_36_61_buffered : std_logic_vector(15 downto 0);
    signal num_blk_62 : std_logic_vector(15 downto 0);
    signal num_left_58 : std_logic_vector(15 downto 0);
    signal ptr_deref_139_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_139_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_139_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_139_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_139_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_77 : std_logic_vector(15 downto 0);
    signal type_cast_125_wire : std_logic_vector(15 downto 0);
    signal type_cast_249_wire : std_logic_vector(31 downto 0);
    signal type_cast_267_wire : std_logic_vector(1 downto 0);
    signal type_cast_276_wire : std_logic_vector(63 downto 0);
    signal type_cast_51_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_56_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_66_wire : std_logic_vector(15 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_81_wire_constant : std_logic_vector(15 downto 0);
    signal w1_144 : std_logic_vector(15 downto 0);
    signal w2_148 : std_logic_vector(15 downto 0);
    signal w3_152 : std_logic_vector(15 downto 0);
    signal w4_156 : std_logic_vector(15 downto 0);
    signal winr_67 : std_logic_vector(15 downto 0);
    signal winr_done_194 : std_logic_vector(0 downto 0);
    signal word_read_140 : std_logic_vector(63 downto 0);
    signal word_start_52 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_134_constant_part_of_offset <= "00000000000000";
    array_obj_ref_134_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_134_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_134_resized_base_address <= "00000000000000";
    konst_103_wire_constant <= "00";
    konst_106_wire_constant <= "0000000000000010";
    konst_110_wire_constant <= "01";
    konst_113_wire_constant <= "0000000000000001";
    konst_117_wire_constant <= "10";
    konst_127_wire_constant <= "0000000000000011";
    konst_203_wire_constant <= "0000000000000000";
    konst_205_wire_constant <= "0000000000000001";
    konst_216_wire_constant <= "0000000000000000";
    konst_218_wire_constant <= "0000000000000001";
    konst_231_wire_constant <= "0000000000000001";
    konst_260_wire_constant <= "00000000000000000000000000000011";
    konst_268_wire_constant <= "00";
    konst_274_wire_constant <= "00000000000000000000000000000010";
    konst_278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_295_wire_constant <= "0000000000000100";
    konst_297_wire_constant <= "0000000000000100";
    konst_303_wire_constant <= "0000000000000100";
    konst_306_wire_constant <= "0000000000000100";
    konst_39_wire_constant <= "0000000000000100";
    konst_42_wire_constant <= "0000000000000100";
    konst_85_wire_constant <= "00";
    konst_90_wire_constant <= "00";
    konst_93_wire_constant <= "0000000000000001";
    konst_97_wire_constant <= "01";
    ptr_deref_139_word_offset_0 <= "00000000000000";
    type_cast_51_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_56_wire_constant <= "00";
    type_cast_70_wire_constant <= "0000000000000000";
    type_cast_76_wire_constant <= "0000000000000000";
    type_cast_81_wire_constant <= "0000000000000000";
    phi_stmt_47: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address_281_49_buffered & type_cast_51_wire_constant;
      req <= phi_stmt_47_req_0 & phi_stmt_47_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_47",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_47_ack_0,
          idata => idata,
          odata => address_47,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_47
    phi_stmt_52: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_56_wire_constant & n_word_start_270_57_buffered;
      req <= phi_stmt_52_req_0 & phi_stmt_52_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_52",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_52_ack_0,
          idata => idata,
          odata => word_start_52,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_52
    phi_stmt_58: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_left_289_60_buffered & nl_start_36_61_buffered;
      req <= phi_stmt_58_req_0 & phi_stmt_58_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_58",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_58_ack_0,
          idata => idata,
          odata => num_left_58,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_58
    phi_stmt_62: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_blk_309_64_buffered & type_cast_66_wire;
      req <= phi_stmt_62_req_0 & phi_stmt_62_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_62",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_62_ack_0,
          idata => idata,
          odata => num_blk_62,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_62
    phi_stmt_67: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_70_wire_constant & n_winr_210_71_buffered;
      req <= phi_stmt_67_req_0 & phi_stmt_67_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_67",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_67_ack_0,
          idata => idata,
          odata => winr_67,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_67
    phi_stmt_72: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_col_223_74_buffered & type_cast_76_wire_constant;
      req <= phi_stmt_72_req_0 & phi_stmt_72_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_72",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_72_ack_0,
          idata => idata,
          odata => col_72,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_72
    phi_stmt_77: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row_235_79_buffered & type_cast_81_wire_constant;
      req <= phi_stmt_77_req_0 & phi_stmt_77_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_77",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_77_ack_0,
          idata => idata,
          odata => row_77,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_77
    -- flow-through select operator MUX_207_inst
    MUX_207_wire <= konst_203_wire_constant when (winr_done_194(0) /=  '0') else ADD_u16_u16_206_wire;
    -- flow-through select operator MUX_209_inst
    n_winr_210 <= MUX_207_wire when (flag1_189(0) /=  '0') else winr_67;
    -- flow-through select operator MUX_220_inst
    MUX_220_wire <= konst_216_wire_constant when (col_done_199(0) /=  '0') else ADD_u16_u16_219_wire;
    -- flow-through select operator MUX_222_inst
    n_col_223 <= MUX_220_wire when (AND_u1_u1_214_wire(0) /=  '0') else col_72;
    -- flow-through select operator MUX_234_inst
    n_row_235 <= ADD_u16_u16_232_wire when (AND_u1_u1_229_wire(0) /=  '0') else row_77;
    -- flow-through select operator MUX_269_inst
    n_word_start_270 <= type_cast_267_wire when (flag1_189(0) /=  '0') else konst_268_wire_constant;
    -- flow-through select operator MUX_280_inst
    n_address_281 <= type_cast_276_wire when (flag1_189(0) /=  '0') else ADD_u64_u64_279_wire;
    -- flow-through select operator MUX_288_inst
    n_left_289 <= nl_start_36 when (flag1_189(0) /=  '0') else SUB_u16_u16_287_wire;
    -- flow-through select operator MUX_301_inst
    MUX_301_wire <= SUB_u16_u16_299_wire when (UGT_u16_u1_296_wire(0) /=  '0') else fn_blk_44;
    -- flow-through select operator MUX_307_inst
    MUX_307_wire <= n_left_289 when (ULT_u16_u1_304_wire(0) /=  '0') else konst_306_wire_constant;
    -- flow-through select operator MUX_308_inst
    n_blk_309 <= MUX_301_wire when (flag1_189(0) /=  '0') else MUX_307_wire;
    -- flow-through select operator MUX_43_inst
    fn_blk_44 <= num_cont_buffer when (ULT_u16_u1_40_wire(0) /=  '0') else konst_42_wire_constant;
    slice_143_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_143_inst_req_0;
      slice_143_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_143_inst_req_1;
      slice_143_inst_ack_1<= update_ack(0);
      slice_143_inst: SliceSplitProtocol generic map(name => "slice_143_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w1_144, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_147_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_147_inst_req_0;
      slice_147_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_147_inst_req_1;
      slice_147_inst_ack_1<= update_ack(0);
      slice_147_inst: SliceSplitProtocol generic map(name => "slice_147_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w2_148, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_151_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_151_inst_req_0;
      slice_151_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_151_inst_req_1;
      slice_151_inst_ack_1<= update_ack(0);
      slice_151_inst: SliceSplitProtocol generic map(name => "slice_151_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w3_152, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_155_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_155_inst_req_0;
      slice_155_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_155_inst_req_1;
      slice_155_inst_ack_1<= update_ack(0);
      slice_155_inst: SliceSplitProtocol generic map(name => "slice_155_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w4_156, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_157_delayed_14_0_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_157_delayed_14_0_157_inst_req_0;
      W_c1_157_delayed_14_0_157_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_157_delayed_14_0_157_inst_req_1;
      W_c1_157_delayed_14_0_157_inst_ack_1<= rack(0);
      W_c1_157_delayed_14_0_157_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_157_delayed_14_0_157_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_87,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_157_delayed_14_0_159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_161_delayed_14_0_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_161_delayed_14_0_164_inst_req_0;
      W_c2_161_delayed_14_0_164_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_161_delayed_14_0_164_inst_req_1;
      W_c2_161_delayed_14_0_164_inst_ack_1<= rack(0);
      W_c2_161_delayed_14_0_164_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_161_delayed_14_0_164_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_161_delayed_14_0_166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_165_delayed_14_0_171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_165_delayed_14_0_171_inst_req_0;
      W_c3_165_delayed_14_0_171_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_165_delayed_14_0_171_inst_req_1;
      W_c3_165_delayed_14_0_171_inst_ack_1<= rack(0);
      W_c3_165_delayed_14_0_171_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_165_delayed_14_0_171_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_121,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_165_delayed_14_0_173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_169_delayed_14_0_178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_169_delayed_14_0_178_inst_req_0;
      W_c4_169_delayed_14_0_178_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_169_delayed_14_0_178_inst_req_1;
      W_c4_169_delayed_14_0_178_inst_ack_1<= rack(0);
      W_c4_169_delayed_14_0_178_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_169_delayed_14_0_178_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_169_delayed_14_0_180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_34_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_36 <= tmp_var; -- 
    end process;
    addr_of_135_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_135_final_reg_req_0;
      addr_of_135_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_135_final_reg_req_1;
      addr_of_135_final_reg_ack_1<= rack(0);
      addr_of_135_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_135_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_134_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_281_49_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_281_49_buf_req_0;
      n_address_281_49_buf_ack_0<= wack(0);
      rreq(0) <= n_address_281_49_buf_req_1;
      n_address_281_49_buf_ack_1<= rack(0);
      n_address_281_49_buf : InterlockBuffer generic map ( -- 
        name => "n_address_281_49_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_281_49_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_309_64_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_309_64_buf_req_0;
      n_blk_309_64_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_309_64_buf_req_1;
      n_blk_309_64_buf_ack_1<= rack(0);
      n_blk_309_64_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_309_64_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_309_64_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_223_74_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_223_74_buf_req_0;
      n_col_223_74_buf_ack_0<= wack(0);
      rreq(0) <= n_col_223_74_buf_req_1;
      n_col_223_74_buf_ack_1<= rack(0);
      n_col_223_74_buf : InterlockBuffer generic map ( -- 
        name => "n_col_223_74_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_223_74_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_289_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_289_60_buf_req_0;
      n_left_289_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_289_60_buf_req_1;
      n_left_289_60_buf_ack_1<= rack(0);
      n_left_289_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_289_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_289_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_235_79_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_235_79_buf_req_0;
      n_row_235_79_buf_ack_0<= wack(0);
      rreq(0) <= n_row_235_79_buf_req_1;
      n_row_235_79_buf_ack_1<= rack(0);
      n_row_235_79_buf : InterlockBuffer generic map ( -- 
        name => "n_row_235_79_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_235_79_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_210_71_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_210_71_buf_req_0;
      n_winr_210_71_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_210_71_buf_req_1;
      n_winr_210_71_buf_ack_1<= rack(0);
      n_winr_210_71_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_210_71_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_210_71_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_270_57_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_270_57_buf_req_0;
      n_word_start_270_57_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_270_57_buf_req_1;
      n_word_start_270_57_buf_ack_1<= rack(0);
      n_word_start_270_57_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_270_57_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_270_57_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_36_61_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_36_61_buf_req_0;
      nl_start_36_61_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_36_61_buf_req_1;
      nl_start_36_61_buf_ack_1<= rack(0);
      nl_start_36_61_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_36_61_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_36_61_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_125_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_52(1 downto 0);
      type_cast_125_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_244_inst
    process(MUL_u16_u16_243_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_243_wire(15 downto 0);
      na1_245 <= tmp_var; -- 
    end process;
    -- interlock type_cast_249_inst
    process(n_winr_210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_210(15 downto 0);
      type_cast_249_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_251_inst
    process(MUL_u32_u32_250_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_250_wire(31 downto 0);
      na2_252 <= tmp_var; -- 
    end process;
    -- interlock type_cast_262_inst
    process(AND_u32_u32_261_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_261_wire(15 downto 0);
      na4_263 <= tmp_var; -- 
    end process;
    -- interlock type_cast_267_inst
    process(na4_263) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_263(1 downto 0);
      type_cast_267_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_276_inst
    process(LSHR_u32_u32_275_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_275_wire(31 downto 0);
      type_cast_276_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_32_inst
    process(MUL_u16_u16_31_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_31_wire(15 downto 0);
      m_factor_33 <= tmp_var; -- 
    end process;
    type_cast_66_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_66_inst_req_0;
      type_cast_66_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_66_inst_req_1;
      type_cast_66_inst_ack_1<= rack(0);
      type_cast_66_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_66_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_44,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_66_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_134_index_1_rename
    process(R_address_133_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_133_resized;
      ov(13 downto 0) := iv;
      R_address_133_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_134_index_1_resize
    process(address_47) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_47;
      ov := iv(13 downto 0);
      R_address_133_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_134_root_address_inst
    process(array_obj_ref_134_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_134_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_134_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_addr_0
    process(ptr_deref_139_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_139_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_base_resize
    process(fetch_addr_136) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_136;
      ov := iv(13 downto 0);
      ptr_deref_139_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_gather_scatter
    process(ptr_deref_139_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_data_0;
      ov(63 downto 0) := iv;
      word_read_140 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_root_address_inst
    process(ptr_deref_139_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_139_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_45_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_313_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_45_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_45_branch_req_0,
          ack0 => do_while_stmt_45_branch_ack_0,
          ack1 => do_while_stmt_45_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_126_inst
    process(num_blk_62, type_cast_125_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_62, type_cast_125_wire, tmp_var);
      ADD_u16_u16_126_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_206_inst
    process(winr_67) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_67, konst_205_wire_constant, tmp_var);
      ADD_u16_u16_206_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_219_inst
    process(col_72) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_72, konst_218_wire_constant, tmp_var);
      ADD_u16_u16_219_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_232_inst
    process(row_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_77, konst_231_wire_constant, tmp_var);
      ADD_u16_u16_232_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_242_inst
    process(n_col_223, MUL_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_223, MUL_u16_u16_241_wire, tmp_var);
      ADD_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_294_inst
    process(fn_blk_44, na4_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_44, na4_263, tmp_var);
      ADD_u16_u16_294_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_256_inst
    process(na1_245, na2_252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_245, na2_252, tmp_var);
      na3_257 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_279_inst
    process(address_47) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_47, konst_278_wire_constant, tmp_var);
      ADD_u64_u64_279_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_108_inst
    process(EQ_u2_u1_104_wire, UGT_u16_u1_107_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_104_wire, UGT_u16_u1_107_wire, tmp_var);
      AND_u1_u1_108_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_115_inst
    process(EQ_u2_u1_111_wire, UGT_u16_u1_114_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_111_wire, UGT_u16_u1_114_wire, tmp_var);
      AND_u1_u1_115_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_214_inst
    process(winr_done_194, flag1_189) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_194, flag1_189, tmp_var);
      AND_u1_u1_214_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(col_done_199, flag1_189) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_199, flag1_189, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_229_inst
    process(winr_done_194, AND_u1_u1_228_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_194, AND_u1_u1_228_wire, tmp_var);
      AND_u1_u1_229_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_95_inst
    process(EQ_u2_u1_91_wire, UGT_u16_u1_94_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_91_wire, UGT_u16_u1_94_wire, tmp_var);
      AND_u1_u1_95_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_261_inst
    process(na3_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_257, konst_260_wire_constant, tmp_var);
      AND_u32_u32_261_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_188_inst
    process(num_left_58, num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_58, num_blk_62, tmp_var);
      flag1_189 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_193_inst
    process(winr_67, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_67, rk1_buffer, tmp_var);
      winr_done_194 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_198_inst
    process(col_72, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_72, col1_buffer, tmp_var);
      col_done_199 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_104_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_103_wire_constant, tmp_var);
      EQ_u2_u1_104_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_111_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_110_wire_constant, tmp_var);
      EQ_u2_u1_111_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_118_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_117_wire_constant, tmp_var);
      EQ_u2_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_86_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_85_wire_constant, tmp_var);
      c1_87 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_91_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_90_wire_constant, tmp_var);
      EQ_u2_u1_91_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_98_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_97_wire_constant, tmp_var);
      EQ_u2_u1_98_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_275_inst
    process(na3_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_257, konst_274_wire_constant, tmp_var);
      LSHR_u32_u32_275_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_241_inst
    process(ct_buffer, n_row_235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_235, tmp_var);
      MUL_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_243_inst
    process(chl_in_buffer, ADD_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_242_wire, tmp_var);
      MUL_u16_u16_243_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_31_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_31_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_250_inst
    process(m_factor_33, type_cast_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_33, type_cast_249_wire, tmp_var);
      MUL_u32_u32_250_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_313_inst
    process(n_row_235, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_235, row1_buffer, tmp_var);
      NEQ_u16_u1_313_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_115_wire, EQ_u2_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_115_wire, EQ_u2_u1_118_wire, tmp_var);
      OR_u1_u1_119_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_120_inst
    process(AND_u1_u1_108_wire, OR_u1_u1_119_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_108_wire, OR_u1_u1_119_wire, tmp_var);
      c3_121 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_99_inst
    process(AND_u1_u1_95_wire, EQ_u2_u1_98_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_95_wire, EQ_u2_u1_98_wire, tmp_var);
      c2_100 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_287_inst
    process(num_left_58, num_blk_62) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_58, num_blk_62, tmp_var);
      SUB_u16_u16_287_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_299_inst
    process(konst_297_wire_constant, na4_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_297_wire_constant, na4_263, tmp_var);
      SUB_u16_u16_299_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_107_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_106_wire_constant, tmp_var);
      UGT_u16_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_114_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_113_wire_constant, tmp_var);
      UGT_u16_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_128_inst
    process(ADD_u16_u16_126_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_126_wire, konst_127_wire_constant, tmp_var);
      c4_129 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_296_inst
    process(ADD_u16_u16_294_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_294_wire, konst_295_wire_constant, tmp_var);
      UGT_u16_u1_296_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_94_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_93_wire_constant, tmp_var);
      UGT_u16_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_304_inst
    process(n_left_289) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_289, konst_303_wire_constant, tmp_var);
      ULT_u16_u1_304_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_40_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_39_wire_constant, tmp_var);
      ULT_u16_u1_40_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_134_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_133_scaled;
      array_obj_ref_134_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_134_index_offset_req_0;
      array_obj_ref_134_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_134_index_offset_req_1;
      array_obj_ref_134_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_139_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_139_load_0_req_0;
      ptr_deref_139_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_139_load_0_req_1;
      ptr_deref_139_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_139_word_address_0;
      ptr_deref_139_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_175_inst WPIPE_input_pipe1_168_inst WPIPE_input_pipe1_161_inst WPIPE_input_pipe1_182_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_175_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_168_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_161_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_182_inst_req_0;
      WPIPE_input_pipe1_175_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_168_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_161_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_182_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_175_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_168_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_161_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_182_inst_req_1;
      WPIPE_input_pipe1_175_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_168_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_161_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_182_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_169_delayed_14_0_180(0);
      guard_vector(1)  <= c1_157_delayed_14_0_159(0);
      guard_vector(2)  <= c2_161_delayed_14_0_166(0);
      guard_vector(3)  <= c3_165_delayed_14_0_173(0);
      data_in <= w3_152 & w2_148 & w1_144 & w4_156;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(135 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1129_start: Boolean;
  signal convolution3D_CP_1129_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      pp : in  std_logic_vector(7 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_556_inst_req_0 : boolean;
  signal type_cast_661_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_644_inst_ack_1 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal type_cast_635_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_req_0 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_606_inst_req_0 : boolean;
  signal type_cast_535_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_ack_1 : boolean;
  signal type_cast_548_inst_req_1 : boolean;
  signal type_cast_560_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_ack_0 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal type_cast_548_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_ack_0 : boolean;
  signal type_cast_585_inst_ack_1 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal type_cast_560_inst_ack_1 : boolean;
  signal type_cast_635_inst_ack_1 : boolean;
  signal type_cast_573_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_req_1 : boolean;
  signal type_cast_535_inst_ack_1 : boolean;
  signal array_obj_ref_1091_index_offset_ack_1 : boolean;
  signal type_cast_548_inst_ack_1 : boolean;
  signal type_cast_635_inst_req_1 : boolean;
  signal type_cast_548_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_556_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_ack_0 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal type_cast_648_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_581_inst_ack_1 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_ack_0 : boolean;
  signal type_cast_560_inst_req_0 : boolean;
  signal type_cast_573_inst_req_1 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_581_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_581_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_556_inst_req_1 : boolean;
  signal type_cast_657_inst_ack_1 : boolean;
  signal type_cast_635_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_606_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_ack_1 : boolean;
  signal type_cast_585_inst_req_1 : boolean;
  signal type_cast_1283_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_631_inst_ack_1 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_581_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_644_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_556_inst_ack_0 : boolean;
  signal type_cast_535_inst_req_1 : boolean;
  signal type_cast_535_inst_req_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal type_cast_648_inst_req_1 : boolean;
  signal type_cast_560_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_req_0 : boolean;
  signal type_cast_1301_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_req_1 : boolean;
  signal type_cast_657_inst_req_1 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal type_cast_585_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_ack_0 : boolean;
  signal type_cast_523_inst_req_0 : boolean;
  signal type_cast_523_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_req_1 : boolean;
  signal type_cast_585_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_644_inst_req_0 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal type_cast_677_inst_req_1 : boolean;
  signal type_cast_1102_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_ack_1 : boolean;
  signal if_stmt_685_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_631_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_606_inst_req_1 : boolean;
  signal type_cast_677_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_req_1 : boolean;
  signal type_cast_677_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_644_inst_ack_0 : boolean;
  signal if_stmt_685_branch_req_0 : boolean;
  signal type_cast_657_inst_ack_0 : boolean;
  signal type_cast_1301_inst_ack_0 : boolean;
  signal type_cast_677_inst_ack_0 : boolean;
  signal type_cast_1102_inst_ack_1 : boolean;
  signal type_cast_657_inst_req_0 : boolean;
  signal if_stmt_685_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_req_0 : boolean;
  signal type_cast_705_inst_req_1 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_705_inst_ack_1 : boolean;
  signal type_cast_661_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_ack_0 : boolean;
  signal type_cast_705_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_705_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_631_inst_ack_0 : boolean;
  signal type_cast_1204_inst_ack_0 : boolean;
  signal ptr_deref_1095_store_0_ack_0 : boolean;
  signal array_obj_ref_1091_index_offset_ack_0 : boolean;
  signal array_obj_ref_1091_index_offset_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_631_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_606_inst_ack_0 : boolean;
  signal type_cast_661_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_req_1 : boolean;
  signal type_cast_523_inst_ack_1 : boolean;
  signal type_cast_661_inst_ack_0 : boolean;
  signal type_cast_510_inst_ack_1 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal type_cast_510_inst_req_1 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal addr_of_1245_final_reg_req_0 : boolean;
  signal type_cast_523_inst_req_1 : boolean;
  signal addr_of_1245_final_reg_ack_0 : boolean;
  signal type_cast_1045_inst_req_0 : boolean;
  signal addr_of_1092_final_reg_req_1 : boolean;
  signal type_cast_1045_inst_ack_0 : boolean;
  signal addr_of_1092_final_reg_ack_1 : boolean;
  signal type_cast_1204_inst_req_1 : boolean;
  signal array_obj_ref_1244_index_offset_req_0 : boolean;
  signal array_obj_ref_1244_index_offset_ack_0 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal type_cast_1045_inst_req_1 : boolean;
  signal type_cast_1045_inst_ack_1 : boolean;
  signal ptr_deref_1095_store_0_req_1 : boolean;
  signal array_obj_ref_1244_index_offset_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_456_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_456_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_456_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_456_inst_ack_1 : boolean;
  signal type_cast_460_inst_req_0 : boolean;
  signal type_cast_460_inst_ack_0 : boolean;
  signal type_cast_460_inst_req_1 : boolean;
  signal type_cast_460_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_1 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_481_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_481_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_481_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_481_inst_ack_1 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_ack_1 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal type_cast_498_inst_req_1 : boolean;
  signal type_cast_498_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_506_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_506_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_506_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_506_inst_ack_1 : boolean;
  signal type_cast_510_inst_req_0 : boolean;
  signal type_cast_510_inst_ack_0 : boolean;
  signal type_cast_721_inst_req_0 : boolean;
  signal type_cast_721_inst_ack_0 : boolean;
  signal type_cast_721_inst_req_1 : boolean;
  signal type_cast_721_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_ack_0 : boolean;
  signal type_cast_1204_inst_req_0 : boolean;
  signal ptr_deref_1095_store_0_req_0 : boolean;
  signal type_cast_730_inst_req_0 : boolean;
  signal type_cast_730_inst_ack_0 : boolean;
  signal type_cast_730_inst_req_1 : boolean;
  signal type_cast_730_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_req_0 : boolean;
  signal type_cast_740_inst_req_0 : boolean;
  signal type_cast_740_inst_ack_0 : boolean;
  signal type_cast_1102_inst_ack_0 : boolean;
  signal type_cast_740_inst_req_1 : boolean;
  signal type_cast_740_inst_ack_1 : boolean;
  signal phi_stmt_998_req_0 : boolean;
  signal type_cast_1301_inst_req_0 : boolean;
  signal array_obj_ref_1244_index_offset_ack_1 : boolean;
  signal type_cast_1195_inst_ack_1 : boolean;
  signal type_cast_1195_inst_req_1 : boolean;
  signal type_cast_1102_inst_req_0 : boolean;
  signal array_obj_ref_775_index_offset_req_0 : boolean;
  signal array_obj_ref_775_index_offset_ack_0 : boolean;
  signal array_obj_ref_1091_index_offset_req_0 : boolean;
  signal array_obj_ref_775_index_offset_req_1 : boolean;
  signal if_stmt_1152_branch_ack_0 : boolean;
  signal array_obj_ref_775_index_offset_ack_1 : boolean;
  signal type_cast_1301_inst_req_1 : boolean;
  signal type_cast_1252_inst_ack_1 : boolean;
  signal addr_of_776_final_reg_req_0 : boolean;
  signal if_stmt_1152_branch_ack_1 : boolean;
  signal addr_of_776_final_reg_ack_0 : boolean;
  signal type_cast_1252_inst_req_1 : boolean;
  signal addr_of_776_final_reg_req_1 : boolean;
  signal addr_of_776_final_reg_ack_1 : boolean;
  signal type_cast_1195_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_779_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_779_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_779_inst_req_1 : boolean;
  signal if_stmt_1152_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_779_inst_ack_1 : boolean;
  signal type_cast_1319_inst_req_0 : boolean;
  signal type_cast_1195_inst_req_0 : boolean;
  signal type_cast_783_inst_req_0 : boolean;
  signal type_cast_783_inst_ack_0 : boolean;
  signal type_cast_783_inst_req_1 : boolean;
  signal type_cast_783_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_792_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_req_1 : boolean;
  signal type_cast_1252_inst_ack_0 : boolean;
  signal type_cast_796_inst_req_0 : boolean;
  signal type_cast_796_inst_ack_0 : boolean;
  signal type_cast_1252_inst_req_0 : boolean;
  signal type_cast_796_inst_req_1 : boolean;
  signal type_cast_1114_inst_ack_1 : boolean;
  signal type_cast_796_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_0 : boolean;
  signal type_cast_1114_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1279_inst_req_0 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal type_cast_1114_inst_ack_0 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_req_1 : boolean;
  signal type_cast_1186_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_req_0 : boolean;
  signal type_cast_1114_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_828_inst_ack_1 : boolean;
  signal type_cast_1186_inst_req_1 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal if_stmt_1052_branch_ack_0 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal type_cast_1751_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_1 : boolean;
  signal type_cast_1004_inst_req_0 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal type_cast_850_inst_req_1 : boolean;
  signal type_cast_850_inst_ack_1 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_req_1 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_864_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_req_1 : boolean;
  signal type_cast_1265_inst_ack_1 : boolean;
  signal type_cast_1265_inst_req_1 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal type_cast_868_inst_req_0 : boolean;
  signal type_cast_868_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1248_inst_ack_1 : boolean;
  signal type_cast_868_inst_req_1 : boolean;
  signal type_cast_868_inst_ack_1 : boolean;
  signal type_cast_1751_inst_ack_1 : boolean;
  signal type_cast_1283_inst_ack_1 : boolean;
  signal type_cast_1209_inst_ack_1 : boolean;
  signal type_cast_1209_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_req_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_882_inst_ack_1 : boolean;
  signal type_cast_1265_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1248_inst_req_1 : boolean;
  signal type_cast_886_inst_req_0 : boolean;
  signal type_cast_886_inst_ack_0 : boolean;
  signal type_cast_886_inst_req_1 : boolean;
  signal type_cast_886_inst_ack_1 : boolean;
  signal type_cast_1319_inst_ack_1 : boolean;
  signal type_cast_1283_inst_req_1 : boolean;
  signal type_cast_1209_inst_ack_0 : boolean;
  signal type_cast_1209_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_900_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_900_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_900_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_900_inst_ack_1 : boolean;
  signal type_cast_1177_inst_ack_1 : boolean;
  signal addr_of_1245_final_reg_ack_1 : boolean;
  signal type_cast_904_inst_req_0 : boolean;
  signal type_cast_904_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1248_inst_ack_0 : boolean;
  signal type_cast_904_inst_req_1 : boolean;
  signal type_cast_904_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_ack_0 : boolean;
  signal type_cast_1319_inst_req_1 : boolean;
  signal type_cast_1177_inst_req_1 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_1 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1248_inst_req_0 : boolean;
  signal addr_of_1092_final_reg_ack_0 : boolean;
  signal ptr_deref_912_store_0_req_0 : boolean;
  signal ptr_deref_912_store_0_ack_0 : boolean;
  signal addr_of_1092_final_reg_req_0 : boolean;
  signal ptr_deref_912_store_0_req_1 : boolean;
  signal ptr_deref_912_store_0_ack_1 : boolean;
  signal type_cast_1283_inst_ack_0 : boolean;
  signal type_cast_1319_inst_ack_0 : boolean;
  signal if_stmt_926_branch_req_0 : boolean;
  signal if_stmt_1052_branch_ack_1 : boolean;
  signal if_stmt_926_branch_ack_1 : boolean;
  signal if_stmt_926_branch_ack_0 : boolean;
  signal if_stmt_1052_branch_req_0 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1315_inst_req_0 : boolean;
  signal if_stmt_977_branch_req_0 : boolean;
  signal if_stmt_977_branch_ack_1 : boolean;
  signal ptr_deref_1095_store_0_ack_1 : boolean;
  signal if_stmt_977_branch_ack_0 : boolean;
  signal addr_of_1245_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1261_inst_ack_1 : boolean;
  signal type_cast_1204_inst_ack_1 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1026_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1026_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1026_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1026_inst_ack_1 : boolean;
  signal type_cast_960_inst_req_0 : boolean;
  signal type_cast_1030_inst_req_0 : boolean;
  signal type_cast_1030_inst_ack_0 : boolean;
  signal type_cast_1030_inst_req_1 : boolean;
  signal type_cast_1030_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1333_inst_ack_1 : boolean;
  signal type_cast_1771_inst_ack_0 : boolean;
  signal type_cast_1771_inst_req_0 : boolean;
  signal type_cast_1337_inst_req_0 : boolean;
  signal type_cast_1337_inst_ack_0 : boolean;
  signal type_cast_1337_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1824_inst_ack_1 : boolean;
  signal type_cast_1337_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1809_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1824_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1351_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1809_inst_req_1 : boolean;
  signal type_cast_1355_inst_req_0 : boolean;
  signal type_cast_1355_inst_ack_0 : boolean;
  signal type_cast_1355_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1824_inst_ack_0 : boolean;
  signal type_cast_1355_inst_ack_1 : boolean;
  signal phi_stmt_998_req_1 : boolean;
  signal type_cast_1011_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1809_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1809_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1369_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1824_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1369_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1369_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1369_inst_ack_1 : boolean;
  signal type_cast_1373_inst_req_0 : boolean;
  signal type_cast_1373_inst_ack_0 : boolean;
  signal type_cast_1373_inst_req_1 : boolean;
  signal type_cast_1373_inst_ack_1 : boolean;
  signal type_cast_1004_inst_ack_1 : boolean;
  signal type_cast_1011_inst_req_0 : boolean;
  signal phi_stmt_763_req_1 : boolean;
  signal type_cast_1791_inst_ack_1 : boolean;
  signal phi_stmt_763_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1821_inst_ack_1 : boolean;
  signal type_cast_1791_inst_req_1 : boolean;
  signal ptr_deref_1381_store_0_req_0 : boolean;
  signal ptr_deref_1381_store_0_ack_0 : boolean;
  signal ptr_deref_1381_store_0_req_1 : boolean;
  signal ptr_deref_1381_store_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1806_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1806_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_ack_0 : boolean;
  signal if_stmt_1395_branch_req_0 : boolean;
  signal type_cast_1761_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_req_0 : boolean;
  signal type_cast_1761_inst_req_1 : boolean;
  signal if_stmt_1395_branch_ack_1 : boolean;
  signal if_stmt_1395_branch_ack_0 : boolean;
  signal type_cast_766_inst_ack_1 : boolean;
  signal type_cast_1004_inst_req_1 : boolean;
  signal type_cast_766_inst_req_1 : boolean;
  signal type_cast_1761_inst_ack_0 : boolean;
  signal if_stmt_1446_branch_req_0 : boolean;
  signal type_cast_1761_inst_req_0 : boolean;
  signal if_stmt_1446_branch_ack_1 : boolean;
  signal if_stmt_1446_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1812_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1812_inst_req_1 : boolean;
  signal type_cast_1461_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1821_inst_req_1 : boolean;
  signal type_cast_1461_inst_ack_0 : boolean;
  signal type_cast_1461_inst_req_1 : boolean;
  signal type_cast_1461_inst_ack_1 : boolean;
  signal phi_stmt_1005_req_0 : boolean;
  signal phi_stmt_957_ack_0 : boolean;
  signal phi_stmt_957_req_1 : boolean;
  signal type_cast_766_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1499_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1821_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1499_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1499_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1821_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1499_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1806_inst_ack_0 : boolean;
  signal phi_stmt_957_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1806_inst_req_0 : boolean;
  signal phi_stmt_763_ack_0 : boolean;
  signal type_cast_1503_inst_req_0 : boolean;
  signal type_cast_1503_inst_ack_0 : boolean;
  signal type_cast_1503_inst_req_1 : boolean;
  signal type_cast_1503_inst_ack_1 : boolean;
  signal type_cast_1781_inst_ack_1 : boolean;
  signal type_cast_1004_inst_ack_0 : boolean;
  signal type_cast_960_inst_ack_0 : boolean;
  signal type_cast_1518_inst_req_0 : boolean;
  signal type_cast_1518_inst_ack_0 : boolean;
  signal type_cast_1518_inst_req_1 : boolean;
  signal type_cast_1518_inst_ack_1 : boolean;
  signal type_cast_1781_inst_req_1 : boolean;
  signal if_stmt_1525_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1812_inst_ack_0 : boolean;
  signal if_stmt_1525_branch_ack_1 : boolean;
  signal if_stmt_1525_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1812_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1803_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1803_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1803_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1803_inst_req_0 : boolean;
  signal type_cast_1751_inst_ack_0 : boolean;
  signal type_cast_766_inst_req_0 : boolean;
  signal array_obj_ref_1564_index_offset_req_0 : boolean;
  signal array_obj_ref_1564_index_offset_ack_0 : boolean;
  signal type_cast_1781_inst_ack_0 : boolean;
  signal array_obj_ref_1564_index_offset_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1818_inst_ack_1 : boolean;
  signal array_obj_ref_1564_index_offset_ack_1 : boolean;
  signal type_cast_960_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1818_inst_req_1 : boolean;
  signal type_cast_1781_inst_req_0 : boolean;
  signal type_cast_960_inst_req_1 : boolean;
  signal addr_of_1565_final_reg_req_0 : boolean;
  signal addr_of_1565_final_reg_ack_0 : boolean;
  signal addr_of_1565_final_reg_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1818_inst_ack_0 : boolean;
  signal addr_of_1565_final_reg_ack_1 : boolean;
  signal type_cast_1801_inst_ack_1 : boolean;
  signal type_cast_1801_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1818_inst_req_0 : boolean;
  signal type_cast_1801_inst_ack_0 : boolean;
  signal type_cast_1801_inst_req_0 : boolean;
  signal type_cast_1751_inst_req_0 : boolean;
  signal type_cast_1791_inst_ack_0 : boolean;
  signal type_cast_1791_inst_req_0 : boolean;
  signal ptr_deref_1568_store_0_req_0 : boolean;
  signal ptr_deref_1568_store_0_ack_0 : boolean;
  signal ptr_deref_1568_store_0_req_1 : boolean;
  signal ptr_deref_1568_store_0_ack_1 : boolean;
  signal type_cast_1771_inst_ack_1 : boolean;
  signal call_stmt_1575_call_req_0 : boolean;
  signal call_stmt_1575_call_ack_0 : boolean;
  signal call_stmt_1575_call_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1815_inst_ack_1 : boolean;
  signal call_stmt_1575_call_ack_1 : boolean;
  signal type_cast_1771_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1586_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1586_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1586_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1586_inst_ack_1 : boolean;
  signal type_cast_1615_inst_req_0 : boolean;
  signal type_cast_1615_inst_ack_0 : boolean;
  signal type_cast_1615_inst_req_1 : boolean;
  signal type_cast_1615_inst_ack_1 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal type_cast_1634_inst_req_0 : boolean;
  signal type_cast_1634_inst_ack_0 : boolean;
  signal type_cast_1634_inst_req_1 : boolean;
  signal type_cast_1634_inst_ack_1 : boolean;
  signal type_cast_1663_inst_req_0 : boolean;
  signal type_cast_1663_inst_ack_0 : boolean;
  signal type_cast_1663_inst_req_1 : boolean;
  signal type_cast_1663_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1665_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1665_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1665_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1665_inst_ack_1 : boolean;
  signal type_cast_1670_inst_req_0 : boolean;
  signal type_cast_1670_inst_ack_0 : boolean;
  signal type_cast_1670_inst_req_1 : boolean;
  signal type_cast_1670_inst_ack_1 : boolean;
  signal type_cast_1674_inst_req_0 : boolean;
  signal type_cast_1674_inst_ack_0 : boolean;
  signal type_cast_1674_inst_req_1 : boolean;
  signal type_cast_1674_inst_ack_1 : boolean;
  signal call_stmt_1685_call_req_0 : boolean;
  signal call_stmt_1685_call_ack_0 : boolean;
  signal call_stmt_1685_call_req_1 : boolean;
  signal call_stmt_1685_call_ack_1 : boolean;
  signal call_stmt_1692_call_req_0 : boolean;
  signal call_stmt_1692_call_ack_0 : boolean;
  signal call_stmt_1692_call_req_1 : boolean;
  signal call_stmt_1692_call_ack_1 : boolean;
  signal if_stmt_1704_branch_req_0 : boolean;
  signal if_stmt_1704_branch_ack_1 : boolean;
  signal if_stmt_1704_branch_ack_0 : boolean;
  signal type_cast_1714_inst_req_0 : boolean;
  signal type_cast_1714_inst_ack_0 : boolean;
  signal type_cast_1714_inst_req_1 : boolean;
  signal type_cast_1714_inst_ack_1 : boolean;
  signal call_stmt_1718_call_req_0 : boolean;
  signal call_stmt_1718_call_ack_0 : boolean;
  signal call_stmt_1718_call_req_1 : boolean;
  signal call_stmt_1718_call_ack_1 : boolean;
  signal type_cast_1722_inst_req_0 : boolean;
  signal type_cast_1722_inst_ack_0 : boolean;
  signal type_cast_1722_inst_req_1 : boolean;
  signal type_cast_1722_inst_ack_1 : boolean;
  signal type_cast_1731_inst_req_0 : boolean;
  signal type_cast_1731_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_1 : boolean;
  signal type_cast_1731_inst_ack_1 : boolean;
  signal type_cast_1741_inst_req_0 : boolean;
  signal type_cast_1741_inst_ack_0 : boolean;
  signal type_cast_1741_inst_req_1 : boolean;
  signal type_cast_1741_inst_ack_1 : boolean;
  signal type_cast_1011_inst_req_1 : boolean;
  signal type_cast_1011_inst_ack_1 : boolean;
  signal phi_stmt_1005_req_1 : boolean;
  signal phi_stmt_998_ack_0 : boolean;
  signal phi_stmt_1005_ack_0 : boolean;
  signal type_cast_1062_inst_req_0 : boolean;
  signal type_cast_1062_inst_ack_0 : boolean;
  signal type_cast_1062_inst_req_1 : boolean;
  signal type_cast_1062_inst_ack_1 : boolean;
  signal phi_stmt_1059_req_0 : boolean;
  signal phi_stmt_1059_ack_0 : boolean;
  signal phi_stmt_1232_req_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal phi_stmt_1232_req_1 : boolean;
  signal phi_stmt_1232_ack_0 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal phi_stmt_1426_req_0 : boolean;
  signal phi_stmt_1426_req_1 : boolean;
  signal phi_stmt_1426_ack_0 : boolean;
  signal phi_stmt_1471_req_0 : boolean;
  signal phi_stmt_1478_req_0 : boolean;
  signal type_cast_1477_inst_req_0 : boolean;
  signal type_cast_1477_inst_ack_0 : boolean;
  signal type_cast_1477_inst_req_1 : boolean;
  signal type_cast_1477_inst_ack_1 : boolean;
  signal phi_stmt_1471_req_1 : boolean;
  signal type_cast_1484_inst_req_0 : boolean;
  signal type_cast_1484_inst_ack_0 : boolean;
  signal type_cast_1484_inst_req_1 : boolean;
  signal type_cast_1484_inst_ack_1 : boolean;
  signal phi_stmt_1478_req_1 : boolean;
  signal phi_stmt_1471_ack_0 : boolean;
  signal phi_stmt_1478_ack_0 : boolean;
  signal type_cast_1535_inst_req_0 : boolean;
  signal type_cast_1535_inst_ack_0 : boolean;
  signal type_cast_1535_inst_req_1 : boolean;
  signal type_cast_1535_inst_ack_1 : boolean;
  signal phi_stmt_1532_req_0 : boolean;
  signal phi_stmt_1532_ack_0 : boolean;
  signal phi_stmt_1643_req_1 : boolean;
  signal type_cast_1646_inst_req_0 : boolean;
  signal type_cast_1646_inst_ack_0 : boolean;
  signal type_cast_1646_inst_req_1 : boolean;
  signal type_cast_1646_inst_ack_1 : boolean;
  signal phi_stmt_1643_req_0 : boolean;
  signal phi_stmt_1643_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1129_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1129_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1129_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1129_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1129: Block -- control-path 
    signal convolution3D_CP_1129_elements: BooleanArray(374 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1129_elements(0) <= convolution3D_CP_1129_start;
    convolution3D_CP_1129_symbol <= convolution3D_CP_1129_elements(306);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_453/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/branch_block_stmt_453__entry__
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684__entry__
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_update_start_
      -- CP-element group 0: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Update/$entry
      -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_548_inst_req_1); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_560_inst_req_1); -- 
    cr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_635_inst_req_1); -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_610_inst_req_1); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_573_inst_req_1); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_585_inst_req_1); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_598_inst_req_1); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_535_inst_req_1); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_648_inst_req_1); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_657_inst_req_1); -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_623_inst_req_1); -- 
    cr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_677_inst_req_1); -- 
    cr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_661_inst_req_1); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_510_inst_req_1); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_523_inst_req_1); -- 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => RPIPE_maxpool_input_pipe_456_inst_req_0); -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_460_inst_req_1); -- 
    cr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_473_inst_req_1); -- 
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_485_inst_req_1); -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(0), ack => type_cast_498_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_update_start_
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Update/cr
      -- 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_456_inst_ack_0, ack => convolution3D_CP_1129_elements(1)); -- 
    cr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(1), ack => RPIPE_maxpool_input_pipe_456_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_456_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Sample/rr
      -- 
    ca_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_456_inst_ack_1, ack => convolution3D_CP_1129_elements(2)); -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(2), ack => type_cast_460_inst_req_0); -- 
    rr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(2), ack => RPIPE_maxpool_input_pipe_469_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Sample/ra
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_460_inst_ack_0, ack => convolution3D_CP_1129_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_460_Update/ca
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_460_inst_ack_1, ack => convolution3D_CP_1129_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_update_start_
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Update/cr
      -- 
    ra_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_0, ack => convolution3D_CP_1129_elements(5)); -- 
    cr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(5), ack => RPIPE_maxpool_input_pipe_469_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_469_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Sample/rr
      -- 
    ca_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_1, ack => convolution3D_CP_1129_elements(6)); -- 
    rr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(6), ack => type_cast_473_inst_req_0); -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(6), ack => RPIPE_maxpool_input_pipe_481_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Sample/ra
      -- 
    ra_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => convolution3D_CP_1129_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_473_Update/ca
      -- 
    ca_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => convolution3D_CP_1129_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_update_start_
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Update/cr
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_481_inst_ack_0, ack => convolution3D_CP_1129_elements(9)); -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(9), ack => RPIPE_maxpool_input_pipe_481_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_481_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Sample/rr
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_481_inst_ack_1, ack => convolution3D_CP_1129_elements(10)); -- 
    rr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(10), ack => type_cast_485_inst_req_0); -- 
    rr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(10), ack => RPIPE_maxpool_input_pipe_494_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Sample/ra
      -- 
    ra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => convolution3D_CP_1129_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_485_Update/ca
      -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => convolution3D_CP_1129_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_update_start_
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Update/cr
      -- 
    ra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_494_inst_ack_0, ack => convolution3D_CP_1129_elements(13)); -- 
    cr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(13), ack => RPIPE_maxpool_input_pipe_494_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_494_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Sample/rr
      -- 
    ca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_494_inst_ack_1, ack => convolution3D_CP_1129_elements(14)); -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(14), ack => type_cast_498_inst_req_0); -- 
    rr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(14), ack => RPIPE_maxpool_input_pipe_506_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Sample/ra
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_0, ack => convolution3D_CP_1129_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_498_Update/ca
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_1, ack => convolution3D_CP_1129_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_update_start_
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Update/cr
      -- 
    ra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_506_inst_ack_0, ack => convolution3D_CP_1129_elements(17)); -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(17), ack => RPIPE_maxpool_input_pipe_506_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_506_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Sample/rr
      -- 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_506_inst_ack_1, ack => convolution3D_CP_1129_elements(18)); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(18), ack => type_cast_510_inst_req_0); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(18), ack => RPIPE_maxpool_input_pipe_519_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Sample/ra
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_0, ack => convolution3D_CP_1129_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_510_Update/$exit
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_1, ack => convolution3D_CP_1129_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_update_start_
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Update/cr
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_519_inst_ack_0, ack => convolution3D_CP_1129_elements(21)); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(21), ack => RPIPE_maxpool_input_pipe_519_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_519_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_sample_start_
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_519_inst_ack_1, ack => convolution3D_CP_1129_elements(22)); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(22), ack => type_cast_523_inst_req_0); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(22), ack => RPIPE_maxpool_input_pipe_531_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Sample/ra
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_0, ack => convolution3D_CP_1129_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_523_Update/$exit
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_1, ack => convolution3D_CP_1129_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_update_start_
      -- CP-element group 25: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_sample_completed_
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_531_inst_ack_0, ack => convolution3D_CP_1129_elements(25)); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(25), ack => RPIPE_maxpool_input_pipe_531_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_531_Update/$exit
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_531_inst_ack_1, ack => convolution3D_CP_1129_elements(26)); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(26), ack => type_cast_535_inst_req_0); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(26), ack => RPIPE_maxpool_input_pipe_544_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Sample/$exit
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_535_inst_ack_0, ack => convolution3D_CP_1129_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_535_update_completed_
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_535_inst_ack_1, ack => convolution3D_CP_1129_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_update_start_
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Update/cr
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_544_inst_ack_0, ack => convolution3D_CP_1129_elements(29)); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(29), ack => RPIPE_maxpool_input_pipe_544_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_544_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Sample/$entry
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_544_inst_ack_1, ack => convolution3D_CP_1129_elements(30)); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(30), ack => type_cast_548_inst_req_0); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(30), ack => RPIPE_maxpool_input_pipe_556_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_sample_completed_
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_0, ack => convolution3D_CP_1129_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_548_update_completed_
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_1, ack => convolution3D_CP_1129_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_update_start_
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Sample/$exit
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_556_inst_ack_0, ack => convolution3D_CP_1129_elements(33)); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(33), ack => RPIPE_maxpool_input_pipe_556_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_556_update_completed_
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_556_inst_ack_1, ack => convolution3D_CP_1129_elements(34)); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(34), ack => type_cast_560_inst_req_0); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(34), ack => RPIPE_maxpool_input_pipe_569_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Sample/ra
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_560_inst_ack_0, ack => convolution3D_CP_1129_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_560_Update/ca
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_560_inst_ack_1, ack => convolution3D_CP_1129_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_update_start_
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Update/cr
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_569_inst_ack_0, ack => convolution3D_CP_1129_elements(37)); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(37), ack => RPIPE_maxpool_input_pipe_569_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_569_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_sample_start_
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_569_inst_ack_1, ack => convolution3D_CP_1129_elements(38)); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(38), ack => type_cast_573_inst_req_0); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(38), ack => RPIPE_maxpool_input_pipe_581_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_sample_completed_
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => convolution3D_CP_1129_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_573_update_completed_
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_1, ack => convolution3D_CP_1129_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_update_start_
      -- CP-element group 41: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_sample_completed_
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_581_inst_ack_0, ack => convolution3D_CP_1129_elements(41)); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(41), ack => RPIPE_maxpool_input_pipe_581_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_581_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Sample/$entry
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_581_inst_ack_1, ack => convolution3D_CP_1129_elements(42)); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(42), ack => type_cast_585_inst_req_0); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(42), ack => RPIPE_maxpool_input_pipe_594_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Sample/ra
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_0, ack => convolution3D_CP_1129_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_585_update_completed_
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_1, ack => convolution3D_CP_1129_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_update_start_
      -- CP-element group 45: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_sample_completed_
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_594_inst_ack_0, ack => convolution3D_CP_1129_elements(45)); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(45), ack => RPIPE_maxpool_input_pipe_594_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_594_update_completed_
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_594_inst_ack_1, ack => convolution3D_CP_1129_elements(46)); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(46), ack => type_cast_598_inst_req_0); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(46), ack => RPIPE_maxpool_input_pipe_606_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_sample_completed_
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => convolution3D_CP_1129_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_598_Update/$exit
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => convolution3D_CP_1129_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_update_start_
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_606_inst_ack_0, ack => convolution3D_CP_1129_elements(49)); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(49), ack => RPIPE_maxpool_input_pipe_606_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_606_Update/$exit
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_606_inst_ack_1, ack => convolution3D_CP_1129_elements(50)); -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(50), ack => type_cast_610_inst_req_0); -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(50), ack => RPIPE_maxpool_input_pipe_619_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Sample/ra
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => convolution3D_CP_1129_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_610_update_completed_
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => convolution3D_CP_1129_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_update_start_
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Update/cr
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_619_inst_ack_0, ack => convolution3D_CP_1129_elements(53)); -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(53), ack => RPIPE_maxpool_input_pipe_619_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_619_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Sample/$entry
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_619_inst_ack_1, ack => convolution3D_CP_1129_elements(54)); -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(54), ack => type_cast_623_inst_req_0); -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(54), ack => RPIPE_maxpool_input_pipe_631_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_sample_completed_
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => convolution3D_CP_1129_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_623_update_completed_
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => convolution3D_CP_1129_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_update_start_
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Sample/$exit
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_631_inst_ack_0, ack => convolution3D_CP_1129_elements(57)); -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(57), ack => RPIPE_maxpool_input_pipe_631_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_631_Update/$exit
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_631_inst_ack_1, ack => convolution3D_CP_1129_elements(58)); -- 
    rr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(58), ack => type_cast_635_inst_req_0); -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(58), ack => RPIPE_maxpool_input_pipe_644_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_sample_completed_
      -- 
    ra_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_0, ack => convolution3D_CP_1129_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_635_Update/$exit
      -- 
    ca_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_635_inst_ack_1, ack => convolution3D_CP_1129_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_update_start_
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_644_inst_ack_0, ack => convolution3D_CP_1129_elements(61)); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(61), ack => RPIPE_maxpool_input_pipe_644_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/RPIPE_maxpool_input_pipe_644_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_sample_start_
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_644_inst_ack_1, ack => convolution3D_CP_1129_elements(62)); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(62), ack => type_cast_648_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_0, ack => convolution3D_CP_1129_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_648_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_1, ack => convolution3D_CP_1129_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Sample/$entry
      -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(65), ack => type_cast_657_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(12) & convolution3D_CP_1129_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Sample/$exit
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_657_inst_ack_0, ack => convolution3D_CP_1129_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_657_update_completed_
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_657_inst_ack_1, ack => convolution3D_CP_1129_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_sample_start_
      -- 
    rr_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(68), ack => type_cast_661_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(20) & convolution3D_CP_1129_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Sample/ra
      -- 
    ra_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_0, ack => convolution3D_CP_1129_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_661_Update/$exit
      -- 
    ca_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_1, ack => convolution3D_CP_1129_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Sample/rr
      -- 
    rr_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(71), ack => type_cast_677_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(4) & convolution3D_CP_1129_elements(8) & convolution3D_CP_1129_elements(67) & convolution3D_CP_1129_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_sample_completed_
      -- 
    ra_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_0, ack => convolution3D_CP_1129_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/type_cast_677_Update/$exit
      -- 
    ca_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_677_inst_ack_1, ack => convolution3D_CP_1129_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_453/R_cmp387_686_place
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684__exit__
      -- CP-element group 74: 	 branch_block_stmt_453/if_stmt_685__entry__
      -- CP-element group 74: 	 branch_block_stmt_453/assign_stmt_457_to_assign_stmt_684/$exit
      -- 
    branch_req_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(74), ack => if_stmt_685_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(28) & convolution3D_CP_1129_elements(32) & convolution3D_CP_1129_elements(36) & convolution3D_CP_1129_elements(40) & convolution3D_CP_1129_elements(44) & convolution3D_CP_1129_elements(48) & convolution3D_CP_1129_elements(52) & convolution3D_CP_1129_elements(56) & convolution3D_CP_1129_elements(60) & convolution3D_CP_1129_elements(64) & convolution3D_CP_1129_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_453/if_stmt_685_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_453/if_stmt_685_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_update_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_update_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/entry_bbx_xnph389
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/merge_stmt_691__exit__
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760__entry__
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_update_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_update_start_
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_453/merge_stmt_691_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_453/merge_stmt_691_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_453/merge_stmt_691_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/entry_bbx_xnph389_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_453/entry_bbx_xnph389_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_453/merge_stmt_691_PhiReqMerge
      -- 
    if_choice_transition_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_685_branch_ack_1, ack => convolution3D_CP_1129_elements(75)); -- 
    cr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_705_inst_req_1); -- 
    rr_1757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_705_inst_req_0); -- 
    rr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_721_inst_req_0); -- 
    cr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_721_inst_req_1); -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_730_inst_req_0); -- 
    cr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_730_inst_req_1); -- 
    cr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(75), ack => type_cast_740_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	313 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_453/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_453/if_stmt_685_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_453/if_stmt_685_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/$entry
      -- CP-element group 76: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_685_branch_ack_0, ack => convolution3D_CP_1129_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Sample/ra
      -- 
    ra_1758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_0, ack => convolution3D_CP_1129_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_705_update_completed_
      -- 
    ca_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_705_inst_ack_1, ack => convolution3D_CP_1129_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Sample/ra
      -- 
    ra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_721_inst_ack_0, ack => convolution3D_CP_1129_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_721_Update/ca
      -- 
    ca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_721_inst_ack_1, ack => convolution3D_CP_1129_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Sample/ra
      -- 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_730_inst_ack_0, ack => convolution3D_CP_1129_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_730_Update/ca
      -- 
    ca_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_730_inst_ack_1, ack => convolution3D_CP_1129_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Sample/rr
      -- 
    rr_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(83), ack => type_cast_740_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(80) & convolution3D_CP_1129_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Sample/ra
      -- 
    ra_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_0, ack => convolution3D_CP_1129_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/type_cast_740_Update/ca
      -- 
    ca_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_740_inst_ack_1, ack => convolution3D_CP_1129_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	307 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760/$exit
      -- CP-element group 86: 	 branch_block_stmt_453/assign_stmt_696_to_assign_stmt_760__exit__
      -- CP-element group 86: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/$entry
      -- CP-element group 86: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(78) & convolution3D_CP_1129_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	312 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Sample/ack
      -- 
    ack_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_775_index_offset_ack_0, ack => convolution3D_CP_1129_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	312 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_request/req
      -- 
    ack_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_775_index_offset_ack_1, ack => convolution3D_CP_1129_elements(88)); -- 
    req_1848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(88), ack => addr_of_776_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_request/ack
      -- 
    ack_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_776_final_reg_ack_0, ack => convolution3D_CP_1129_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	312 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_word_addrgen/root_register_ack
      -- 
    ack_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_776_final_reg_ack_1, ack => convolution3D_CP_1129_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	312 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_update_start_
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Update/cr
      -- 
    ra_1863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_779_inst_ack_0, ack => convolution3D_CP_1129_elements(91)); -- 
    cr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(91), ack => RPIPE_maxpool_input_pipe_779_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Sample/rr
      -- 
    ca_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_779_inst_ack_1, ack => convolution3D_CP_1129_elements(92)); -- 
    rr_1876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(92), ack => type_cast_783_inst_req_0); -- 
    rr_1890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(92), ack => RPIPE_maxpool_input_pipe_792_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Sample/ra
      -- 
    ra_1877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_0, ack => convolution3D_CP_1129_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	312 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Update/ca
      -- 
    ca_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_1, ack => convolution3D_CP_1129_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_update_start_
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Update/cr
      -- 
    ra_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_792_inst_ack_0, ack => convolution3D_CP_1129_elements(95)); -- 
    cr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(95), ack => RPIPE_maxpool_input_pipe_792_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_792_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Sample/rr
      -- 
    ca_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_792_inst_ack_1, ack => convolution3D_CP_1129_elements(96)); -- 
    rr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(96), ack => type_cast_796_inst_req_0); -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(96), ack => RPIPE_maxpool_input_pipe_810_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Sample/ra
      -- 
    ra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_0, ack => convolution3D_CP_1129_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	312 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Update/ca
      -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_796_inst_ack_1, ack => convolution3D_CP_1129_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_update_start_
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Update/cr
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_0, ack => convolution3D_CP_1129_elements(99)); -- 
    cr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(99), ack => RPIPE_maxpool_input_pipe_810_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_810_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Sample/rr
      -- 
    ca_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_1, ack => convolution3D_CP_1129_elements(100)); -- 
    rr_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(100), ack => type_cast_814_inst_req_0); -- 
    rr_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(100), ack => RPIPE_maxpool_input_pipe_828_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Sample/ra
      -- 
    ra_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => convolution3D_CP_1129_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	312 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Update/ca
      -- 
    ca_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => convolution3D_CP_1129_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_update_start_
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Update/cr
      -- 
    ra_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_828_inst_ack_0, ack => convolution3D_CP_1129_elements(103)); -- 
    cr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(103), ack => RPIPE_maxpool_input_pipe_828_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_828_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Sample/rr
      -- 
    ca_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_828_inst_ack_1, ack => convolution3D_CP_1129_elements(104)); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(104), ack => type_cast_832_inst_req_0); -- 
    rr_1974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(104), ack => RPIPE_maxpool_input_pipe_846_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Sample/ra
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => convolution3D_CP_1129_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	312 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Update/ca
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => convolution3D_CP_1129_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_update_start_
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Update/cr
      -- 
    ra_1975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_0, ack => convolution3D_CP_1129_elements(107)); -- 
    cr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(107), ack => RPIPE_maxpool_input_pipe_846_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_846_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Sample/rr
      -- 
    ca_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_1, ack => convolution3D_CP_1129_elements(108)); -- 
    rr_1988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(108), ack => type_cast_850_inst_req_0); -- 
    rr_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(108), ack => RPIPE_maxpool_input_pipe_864_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Sample/ra
      -- 
    ra_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => convolution3D_CP_1129_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	312 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Update/ca
      -- 
    ca_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_1, ack => convolution3D_CP_1129_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_update_start_
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Update/cr
      -- 
    ra_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_864_inst_ack_0, ack => convolution3D_CP_1129_elements(111)); -- 
    cr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(111), ack => RPIPE_maxpool_input_pipe_864_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_864_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Sample/rr
      -- 
    ca_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_864_inst_ack_1, ack => convolution3D_CP_1129_elements(112)); -- 
    rr_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(112), ack => type_cast_868_inst_req_0); -- 
    rr_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(112), ack => RPIPE_maxpool_input_pipe_882_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Sample/ra
      -- 
    ra_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_0, ack => convolution3D_CP_1129_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	312 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Update/ca
      -- 
    ca_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_1, ack => convolution3D_CP_1129_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_update_start_
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Update/cr
      -- 
    ra_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_882_inst_ack_0, ack => convolution3D_CP_1129_elements(115)); -- 
    cr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(115), ack => RPIPE_maxpool_input_pipe_882_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_882_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Sample/rr
      -- 
    ca_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_882_inst_ack_1, ack => convolution3D_CP_1129_elements(116)); -- 
    rr_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(116), ack => type_cast_886_inst_req_0); -- 
    rr_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(116), ack => RPIPE_maxpool_input_pipe_900_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Sample/ra
      -- 
    ra_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_886_inst_ack_0, ack => convolution3D_CP_1129_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	312 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Update/ca
      -- 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_886_inst_ack_1, ack => convolution3D_CP_1129_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_update_start_
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Update/cr
      -- 
    ra_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_900_inst_ack_0, ack => convolution3D_CP_1129_elements(119)); -- 
    cr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(119), ack => RPIPE_maxpool_input_pipe_900_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_900_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Sample/rr
      -- 
    ca_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_900_inst_ack_1, ack => convolution3D_CP_1129_elements(120)); -- 
    rr_2072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(120), ack => type_cast_904_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Sample/ra
      -- 
    ra_2073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_0, ack => convolution3D_CP_1129_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	312 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Update/ca
      -- 
    ca_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_904_inst_ack_1, ack => convolution3D_CP_1129_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/ptr_deref_912_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/ptr_deref_912_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/ptr_deref_912_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/ptr_deref_912_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/word_0/rr
      -- 
    rr_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(123), ack => ptr_deref_912_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(90) & convolution3D_CP_1129_elements(94) & convolution3D_CP_1129_elements(98) & convolution3D_CP_1129_elements(102) & convolution3D_CP_1129_elements(106) & convolution3D_CP_1129_elements(110) & convolution3D_CP_1129_elements(114) & convolution3D_CP_1129_elements(118) & convolution3D_CP_1129_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Sample/word_access_start/word_0/ra
      -- 
    ra_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_912_store_0_ack_0, ack => convolution3D_CP_1129_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	312 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/word_0/ca
      -- 
    ca_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_912_store_0_ack_1, ack => convolution3D_CP_1129_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925__exit__
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926__entry__
      -- CP-element group 126: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/$exit
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_453/R_exitcond33_927_place
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_453/if_stmt_926_else_link/$entry
      -- 
    branch_req_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(126), ack => if_stmt_926_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(87) & convolution3D_CP_1129_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	314 
    -- CP-element group 127: 	315 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_453/merge_stmt_932__exit__
      -- CP-element group 127: 	 branch_block_stmt_453/assign_stmt_939_to_assign_stmt_954__entry__
      -- CP-element group 127: 	 branch_block_stmt_453/assign_stmt_939_to_assign_stmt_954__exit__
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_453/merge_stmt_932_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/if_stmt_926_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_453/if_stmt_926_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_453/assign_stmt_939_to_assign_stmt_954/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/assign_stmt_939_to_assign_stmt_954/$exit
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/merge_stmt_932_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_453/merge_stmt_932_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Update/cr
      -- CP-element group 127: 	 branch_block_stmt_453/merge_stmt_932_PhiAck/dummy
      -- 
    if_choice_transition_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_926_branch_ack_1, ack => convolution3D_CP_1129_elements(127)); -- 
    rr_3614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(127), ack => type_cast_960_inst_req_0); -- 
    cr_3619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(127), ack => type_cast_960_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	308 
    -- CP-element group 128: 	309 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/if_stmt_926_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_453/if_stmt_926_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_926_branch_ack_0, ack => convolution3D_CP_1129_elements(128)); -- 
    cr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(128), ack => type_cast_766_inst_req_1); -- 
    rr_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(128), ack => type_cast_766_inst_req_0); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	318 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	337 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_453/if_stmt_977_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_453/if_stmt_977_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_453/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_453/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_453/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_977_branch_ack_1, ack => convolution3D_CP_1129_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	318 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	319 
    -- CP-element group 130: 	320 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_453/merge_stmt_983__exit__
      -- CP-element group 130: 	 branch_block_stmt_453/assign_stmt_989_to_assign_stmt_995__entry__
      -- CP-element group 130: 	 branch_block_stmt_453/assign_stmt_989_to_assign_stmt_995__exit__
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/if_stmt_977_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_453/if_stmt_977_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_453/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_453/assign_stmt_989_to_assign_stmt_995/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/assign_stmt_989_to_assign_stmt_995/$exit
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/merge_stmt_983_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_453/merge_stmt_983_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_453/merge_stmt_983_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_453/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_453/merge_stmt_983_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_453/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- 
    else_choice_transition_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_977_branch_ack_0, ack => convolution3D_CP_1129_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	332 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_update_start_
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Update/cr
      -- 
    ra_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1026_inst_ack_0, ack => convolution3D_CP_1129_elements(131)); -- 
    cr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(131), ack => RPIPE_maxpool_input_pipe_1026_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Sample/rr
      -- 
    ca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1026_inst_ack_1, ack => convolution3D_CP_1129_elements(132)); -- 
    rr_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(132), ack => type_cast_1030_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Sample/ra
      -- 
    ra_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_0, ack => convolution3D_CP_1129_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	332 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Update/ca
      -- 
    ca_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_1, ack => convolution3D_CP_1129_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	332 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Sample/ra
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_0, ack => convolution3D_CP_1129_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	332 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Update/ca
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1045_inst_ack_1, ack => convolution3D_CP_1129_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051__exit__
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052__entry__
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_453/R_cmpx_xi_1053_place
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_else_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_453/if_stmt_1052_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/$exit
      -- 
    branch_req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(137), ack => if_stmt_1052_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(134) & convolution3D_CP_1129_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	322 
    -- CP-element group 138: 	323 
    -- CP-element group 138: 	325 
    -- CP-element group 138: 	326 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/if_stmt_1052_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_453/if_stmt_1052_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1052_branch_ack_1, ack => convolution3D_CP_1129_elements(138)); -- 
    rr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1004_inst_req_0); -- 
    rr_3699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1011_inst_req_0); -- 
    cr_3681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1004_inst_req_1); -- 
    cr_3704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(138), ack => type_cast_1011_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	333 
    -- CP-element group 139: 	334 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_453/if_stmt_1052_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_453/if_stmt_1052_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1052_branch_ack_0, ack => convolution3D_CP_1129_elements(139)); -- 
    rr_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(139), ack => type_cast_1062_inst_req_0); -- 
    cr_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(139), ack => type_cast_1062_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	336 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_sample_complete
      -- 
    ack_2268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_index_offset_ack_0, ack => convolution3D_CP_1129_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	336 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_request/req
      -- CP-element group 141: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_request/$entry
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1091_index_offset_ack_1, ack => convolution3D_CP_1129_elements(141)); -- 
    req_2282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(141), ack => addr_of_1092_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_request/ack
      -- CP-element group 142: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_request/$exit
      -- 
    ack_2283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1092_final_reg_ack_0, ack => convolution3D_CP_1129_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	336 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/word_0/rr
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/ptr_deref_1095_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/ptr_deref_1095_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/ptr_deref_1095_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/ptr_deref_1095_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_base_address_calculated
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1092_final_reg_ack_1, ack => convolution3D_CP_1129_elements(143)); -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(143), ack => ptr_deref_1095_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Sample/$exit
      -- 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1095_store_0_ack_0, ack => convolution3D_CP_1129_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	336 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/word_0/ca
      -- 
    ca_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1095_store_0_ack_1, ack => convolution3D_CP_1129_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	337 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097__exit__
      -- CP-element group 146: 	 branch_block_stmt_453/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/$exit
      -- CP-element group 146: 	 branch_block_stmt_453/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_453/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(140) & convolution3D_CP_1129_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	337 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_sample_completed_
      -- 
    ra_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_0, ack => convolution3D_CP_1129_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	337 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	155 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_update_completed_
      -- 
    ca_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_1, ack => convolution3D_CP_1129_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	337 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Sample/$exit
      -- 
    ra_2364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => convolution3D_CP_1129_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	337 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Update/$exit
      -- 
    ca_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => convolution3D_CP_1129_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	337 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_sample_completed_
      -- 
    ra_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => convolution3D_CP_1129_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	337 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_update_completed_
      -- 
    ca_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => convolution3D_CP_1129_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	337 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_sample_completed_
      -- 
    ra_2392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1114_inst_ack_0, ack => convolution3D_CP_1129_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	337 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_update_completed_
      -- 
    ca_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1114_inst_ack_1, ack => convolution3D_CP_1129_elements(154)); -- 
    -- CP-element group 155:  branch  join  transition  place  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	148 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (10) 
      -- CP-element group 155: 	 branch_block_stmt_453/R_cmp161383_1153_place
      -- CP-element group 155: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151__exit__
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152__entry__
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_else_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_453/if_stmt_1152_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/$exit
      -- 
    branch_req_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(155), ack => if_stmt_1152_branch_req_0); -- 
    convolution3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(148) & convolution3D_CP_1129_elements(150) & convolution3D_CP_1129_elements(152) & convolution3D_CP_1129_elements(154);
      gj_convolution3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	159 
    -- CP-element group 156: 	160 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	162 
    -- CP-element group 156: 	163 
    -- CP-element group 156: 	164 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	168 
    -- CP-element group 156: 	170 
    -- CP-element group 156:  members (42) 
      -- CP-element group 156: 	 branch_block_stmt_453/ifx_xend_bbx_xnph
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_453/merge_stmt_1158__exit__
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229__entry__
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/if_stmt_1152_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_453/if_stmt_1152_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_453/merge_stmt_1158_PhiReqMerge
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_update_start_
      -- CP-element group 156: 	 branch_block_stmt_453/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 156: 	 branch_block_stmt_453/merge_stmt_1158_PhiAck/$entry
      -- CP-element group 156: 	 branch_block_stmt_453/merge_stmt_1158_PhiAck/$exit
      -- CP-element group 156: 	 branch_block_stmt_453/merge_stmt_1158_PhiAck/dummy
      -- 
    if_choice_transition_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_1, ack => convolution3D_CP_1129_elements(156)); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1173_inst_req_1); -- 
    rr_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1173_inst_req_0); -- 
    cr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1204_inst_req_1); -- 
    cr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1195_inst_req_1); -- 
    rr_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1195_inst_req_0); -- 
    cr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1186_inst_req_1); -- 
    rr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1186_inst_req_0); -- 
    cr_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1209_inst_req_1); -- 
    cr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1177_inst_req_1); -- 
    rr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(156), ack => type_cast_1177_inst_req_0); -- 
    -- CP-element group 157:  transition  place  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	347 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_453/ifx_xend_forx_xend215
      -- CP-element group 157: 	 branch_block_stmt_453/if_stmt_1152_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_453/if_stmt_1152_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 157: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/$entry
      -- CP-element group 157: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$entry
      -- 
    else_choice_transition_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1152_branch_ack_0, ack => convolution3D_CP_1129_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_sample_completed_
      -- 
    ra_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convolution3D_CP_1129_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	166 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1173_update_completed_
      -- 
    ca_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convolution3D_CP_1129_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_sample_completed_
      -- 
    ra_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => convolution3D_CP_1129_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1177_update_completed_
      -- 
    ca_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_1, ack => convolution3D_CP_1129_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	156 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_sample_completed_
      -- 
    ra_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_0, ack => convolution3D_CP_1129_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1186_update_completed_
      -- 
    ca_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_1, ack => convolution3D_CP_1129_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_sample_completed_
      -- 
    ra_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1195_inst_ack_0, ack => convolution3D_CP_1129_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1195_update_completed_
      -- 
    ca_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1195_inst_ack_1, ack => convolution3D_CP_1129_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_sample_start_
      -- 
    rr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(166), ack => type_cast_1204_inst_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(159) & convolution3D_CP_1129_elements(161) & convolution3D_CP_1129_elements(163) & convolution3D_CP_1129_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_sample_completed_
      -- 
    ra_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1204_inst_ack_0, ack => convolution3D_CP_1129_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	156 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1204_Update/ca
      -- 
    ca_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1204_inst_ack_1, ack => convolution3D_CP_1129_elements(168)); -- 
    rr_2497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(168), ack => type_cast_1209_inst_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Sample/ra
      -- CP-element group 169: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_sample_completed_
      -- 
    ra_2498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_0, ack => convolution3D_CP_1129_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	156 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	338 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229__exit__
      -- CP-element group 170: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163
      -- CP-element group 170: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/$exit
      -- CP-element group 170: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_453/assign_stmt_1164_to_assign_stmt_1229/type_cast_1209_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/$entry
      -- CP-element group 170: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/$entry
      -- 
    ca_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1209_inst_ack_1, ack => convolution3D_CP_1129_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	343 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Sample/ack
      -- CP-element group 171: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_sample_complete
      -- 
    ack_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1244_index_offset_ack_0, ack => convolution3D_CP_1129_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	343 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_request/req
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_sample_start_
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1244_index_offset_ack_1, ack => convolution3D_CP_1129_elements(172)); -- 
    req_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(172), ack => addr_of_1245_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_request/ack
      -- CP-element group 173: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_sample_completed_
      -- 
    ack_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1245_final_reg_ack_0, ack => convolution3D_CP_1129_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	343 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_word_addrgen/root_register_ack
      -- 
    ack_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1245_final_reg_ack_1, ack => convolution3D_CP_1129_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	343 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_update_start_
      -- CP-element group 175: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_sample_completed_
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1248_inst_ack_0, ack => convolution3D_CP_1129_elements(175)); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(175), ack => RPIPE_maxpool_input_pipe_1248_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_update_completed_
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1248_inst_ack_1, ack => convolution3D_CP_1129_elements(176)); -- 
    rr_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(176), ack => type_cast_1252_inst_req_0); -- 
    rr_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(176), ack => RPIPE_maxpool_input_pipe_1261_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_sample_completed_
      -- 
    ra_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1252_inst_ack_0, ack => convolution3D_CP_1129_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	343 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_update_completed_
      -- 
    ca_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1252_inst_ack_1, ack => convolution3D_CP_1129_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_update_start_
      -- CP-element group 179: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_sample_completed_
      -- 
    ra_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1261_inst_ack_0, ack => convolution3D_CP_1129_elements(179)); -- 
    cr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(179), ack => RPIPE_maxpool_input_pipe_1261_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1261_Update/ca
      -- 
    ca_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1261_inst_ack_1, ack => convolution3D_CP_1129_elements(180)); -- 
    rr_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(180), ack => type_cast_1265_inst_req_0); -- 
    rr_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(180), ack => RPIPE_maxpool_input_pipe_1279_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_sample_completed_
      -- 
    ra_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_0, ack => convolution3D_CP_1129_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	343 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_update_completed_
      -- 
    ca_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_1, ack => convolution3D_CP_1129_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_update_start_
      -- CP-element group 183: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_sample_completed_
      -- 
    ra_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1279_inst_ack_0, ack => convolution3D_CP_1129_elements(183)); -- 
    cr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(183), ack => RPIPE_maxpool_input_pipe_1279_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1279_update_completed_
      -- 
    ca_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1279_inst_ack_1, ack => convolution3D_CP_1129_elements(184)); -- 
    rr_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(184), ack => type_cast_1283_inst_req_0); -- 
    rr_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(184), ack => RPIPE_maxpool_input_pipe_1297_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Sample/ra
      -- 
    ra_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_0, ack => convolution3D_CP_1129_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	343 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Update/$exit
      -- 
    ca_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1283_inst_ack_1, ack => convolution3D_CP_1129_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_update_start_
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Update/cr
      -- 
    ra_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_0, ack => convolution3D_CP_1129_elements(187)); -- 
    cr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(187), ack => RPIPE_maxpool_input_pipe_1297_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1297_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Sample/rr
      -- 
    ca_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_1, ack => convolution3D_CP_1129_elements(188)); -- 
    rr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(188), ack => type_cast_1301_inst_req_0); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(188), ack => RPIPE_maxpool_input_pipe_1315_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_sample_completed_
      -- 
    ra_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_0, ack => convolution3D_CP_1129_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	343 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_update_completed_
      -- 
    ca_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_1, ack => convolution3D_CP_1129_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_update_start_
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Sample/ra
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1315_inst_ack_0, ack => convolution3D_CP_1129_elements(191)); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(191), ack => RPIPE_maxpool_input_pipe_1315_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1315_Update/$exit
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1315_inst_ack_1, ack => convolution3D_CP_1129_elements(192)); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(192), ack => type_cast_1319_inst_req_0); -- 
    rr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(192), ack => RPIPE_maxpool_input_pipe_1333_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Sample/ra
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_0, ack => convolution3D_CP_1129_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	343 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_update_completed_
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1319_inst_ack_1, ack => convolution3D_CP_1129_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_update_start_
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Update/cr
      -- 
    ra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1333_inst_ack_0, ack => convolution3D_CP_1129_elements(195)); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(195), ack => RPIPE_maxpool_input_pipe_1333_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1333_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Sample/rr
      -- 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1333_inst_ack_1, ack => convolution3D_CP_1129_elements(196)); -- 
    rr_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(196), ack => type_cast_1337_inst_req_0); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(196), ack => RPIPE_maxpool_input_pipe_1351_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Sample/ra
      -- 
    ra_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_0, ack => convolution3D_CP_1129_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	343 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Update/ca
      -- 
    ca_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1337_inst_ack_1, ack => convolution3D_CP_1129_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_update_start_
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Update/cr
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1351_inst_ack_0, ack => convolution3D_CP_1129_elements(199)); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(199), ack => RPIPE_maxpool_input_pipe_1351_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1351_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Sample/rr
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1351_inst_ack_1, ack => convolution3D_CP_1129_elements(200)); -- 
    rr_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(200), ack => type_cast_1355_inst_req_0); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(200), ack => RPIPE_maxpool_input_pipe_1369_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Sample/ra
      -- 
    ra_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_0, ack => convolution3D_CP_1129_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	343 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Update/ca
      -- 
    ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1355_inst_ack_1, ack => convolution3D_CP_1129_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_update_start_
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Update/cr
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1369_inst_ack_0, ack => convolution3D_CP_1129_elements(203)); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(203), ack => RPIPE_maxpool_input_pipe_1369_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1369_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Sample/rr
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1369_inst_ack_1, ack => convolution3D_CP_1129_elements(204)); -- 
    rr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(204), ack => type_cast_1373_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Sample/ra
      -- 
    ra_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1373_inst_ack_0, ack => convolution3D_CP_1129_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	343 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Update/ca
      -- 
    ca_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1373_inst_ack_1, ack => convolution3D_CP_1129_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/ptr_deref_1381_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/ptr_deref_1381_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/ptr_deref_1381_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/ptr_deref_1381_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/word_0/rr
      -- 
    rr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(207), ack => ptr_deref_1381_store_0_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(174) & convolution3D_CP_1129_elements(178) & convolution3D_CP_1129_elements(182) & convolution3D_CP_1129_elements(186) & convolution3D_CP_1129_elements(190) & convolution3D_CP_1129_elements(194) & convolution3D_CP_1129_elements(198) & convolution3D_CP_1129_elements(202) & convolution3D_CP_1129_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Sample/word_access_start/word_0/ra
      -- 
    ra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1381_store_0_ack_0, ack => convolution3D_CP_1129_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	343 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/word_0/ca
      -- 
    ca_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1381_store_0_ack_1, ack => convolution3D_CP_1129_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394__exit__
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395__entry__
      -- CP-element group 210: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/$exit
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_453/R_exitcond_1396_place
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_453/if_stmt_1395_else_link/$entry
      -- 
    branch_req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(210), ack => if_stmt_1395_branch_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(171) & convolution3D_CP_1129_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	344 
    -- CP-element group 211: 	345 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_453/merge_stmt_1401_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_453/merge_stmt_1401__exit__
      -- CP-element group 211: 	 branch_block_stmt_453/assign_stmt_1408_to_assign_stmt_1423__entry__
      -- CP-element group 211: 	 branch_block_stmt_453/assign_stmt_1408_to_assign_stmt_1423__exit__
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 211: 	 branch_block_stmt_453/if_stmt_1395_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_453/if_stmt_1395_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 211: 	 branch_block_stmt_453/assign_stmt_1408_to_assign_stmt_1423/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/assign_stmt_1408_to_assign_stmt_1423/$exit
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_453/merge_stmt_1401_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/merge_stmt_1401_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_453/merge_stmt_1401_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1395_branch_ack_1, ack => convolution3D_CP_1129_elements(211)); -- 
    rr_3843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(211), ack => type_cast_1429_inst_req_0); -- 
    cr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(211), ack => type_cast_1429_inst_req_1); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	339 
    -- CP-element group 212: 	340 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_453/if_stmt_1395_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_453/if_stmt_1395_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1395_branch_ack_0, ack => convolution3D_CP_1129_elements(212)); -- 
    rr_3800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(212), ack => type_cast_1238_inst_req_0); -- 
    cr_3805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(212), ack => type_cast_1238_inst_req_1); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	349 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	368 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_453/if_stmt_1446_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_453/if_stmt_1446_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_453/forx_xend215_ifx_xend227
      -- CP-element group 213: 	 branch_block_stmt_453/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_453/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1446_branch_ack_1, ack => convolution3D_CP_1129_elements(213)); -- 
    -- CP-element group 214:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	349 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (18) 
      -- CP-element group 214: 	 branch_block_stmt_453/merge_stmt_1452__exit__
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468__entry__
      -- CP-element group 214: 	 branch_block_stmt_453/if_stmt_1446_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_453/if_stmt_1446_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_453/forx_xend215_bbx_xnphx_xi360
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/$entry
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_update_start_
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_453/forx_xend215_bbx_xnphx_xi360_PhiReq/$entry
      -- CP-element group 214: 	 branch_block_stmt_453/forx_xend215_bbx_xnphx_xi360_PhiReq/$exit
      -- CP-element group 214: 	 branch_block_stmt_453/merge_stmt_1452_PhiReqMerge
      -- CP-element group 214: 	 branch_block_stmt_453/merge_stmt_1452_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_453/merge_stmt_1452_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_453/merge_stmt_1452_PhiAck/dummy
      -- 
    else_choice_transition_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1446_branch_ack_0, ack => convolution3D_CP_1129_elements(214)); -- 
    rr_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(214), ack => type_cast_1461_inst_req_0); -- 
    cr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(214), ack => type_cast_1461_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Sample/ra
      -- 
    ra_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1461_inst_ack_0, ack => convolution3D_CP_1129_elements(215)); -- 
    -- CP-element group 216:  fork  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	350 
    -- CP-element group 216: 	351 
    -- CP-element group 216:  members (11) 
      -- CP-element group 216: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468__exit__
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369
      -- CP-element group 216: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/$exit
      -- CP-element group 216: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_453/assign_stmt_1458_to_assign_stmt_1468/type_cast_1461_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/$entry
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/$entry
      -- CP-element group 216: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/$entry
      -- 
    ca_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1461_inst_ack_1, ack => convolution3D_CP_1129_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	363 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_update_start_
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Update/cr
      -- 
    ra_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1499_inst_ack_0, ack => convolution3D_CP_1129_elements(217)); -- 
    cr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(217), ack => RPIPE_maxpool_input_pipe_1499_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Sample/rr
      -- 
    ca_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1499_inst_ack_1, ack => convolution3D_CP_1129_elements(218)); -- 
    rr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(218), ack => type_cast_1503_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Sample/ra
      -- 
    ra_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1503_inst_ack_0, ack => convolution3D_CP_1129_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	363 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Update/ca
      -- 
    ca_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1503_inst_ack_1, ack => convolution3D_CP_1129_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	363 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Sample/ra
      -- 
    ra_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_0, ack => convolution3D_CP_1129_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	363 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Update/ca
      -- 
    ca_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1518_inst_ack_1, ack => convolution3D_CP_1129_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524__exit__
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525__entry__
      -- CP-element group 223: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/$exit
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_453/R_cmpx_xi368_1526_place
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_453/if_stmt_1525_else_link/$entry
      -- 
    branch_req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(223), ack => if_stmt_1525_branch_req_0); -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(220) & convolution3D_CP_1129_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	353 
    -- CP-element group 224: 	354 
    -- CP-element group 224: 	356 
    -- CP-element group 224: 	357 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_453/if_stmt_1525_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_453/if_stmt_1525_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1525_branch_ack_1, ack => convolution3D_CP_1129_elements(224)); -- 
    rr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1477_inst_req_0); -- 
    cr_3921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1477_inst_req_1); -- 
    rr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1484_inst_req_0); -- 
    cr_3944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(224), ack => type_cast_1484_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	364 
    -- CP-element group 225: 	365 
    -- CP-element group 225:  members (12) 
      -- CP-element group 225: 	 branch_block_stmt_453/if_stmt_1525_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_453/if_stmt_1525_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1525_branch_ack_0, ack => convolution3D_CP_1129_elements(225)); -- 
    rr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(225), ack => type_cast_1535_inst_req_0); -- 
    cr_3980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(225), ack => type_cast_1535_inst_req_1); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	367 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	232 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_sample_complete
      -- CP-element group 226: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Sample/ack
      -- 
    ack_2980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1564_index_offset_ack_0, ack => convolution3D_CP_1129_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	367 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (11) 
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_offset_calculated
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Update/ack
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_request/$entry
      -- CP-element group 227: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_request/req
      -- 
    ack_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1564_index_offset_ack_1, ack => convolution3D_CP_1129_elements(227)); -- 
    req_2994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(227), ack => addr_of_1565_final_reg_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_request/$exit
      -- CP-element group 228: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_request/ack
      -- 
    ack_2995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1565_final_reg_ack_0, ack => convolution3D_CP_1129_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	367 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (28) 
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_complete/ack
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/ptr_deref_1568_Split/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/ptr_deref_1568_Split/$exit
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/ptr_deref_1568_Split/split_req
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/ptr_deref_1568_Split/split_ack
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/word_0/rr
      -- 
    ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1565_final_reg_ack_1, ack => convolution3D_CP_1129_elements(229)); -- 
    rr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(229), ack => ptr_deref_1568_store_0_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Sample/word_access_start/word_0/ra
      -- 
    ra_3039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1568_store_0_ack_0, ack => convolution3D_CP_1129_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	367 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/word_0/ca
      -- 
    ca_3050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1568_store_0_ack_1, ack => convolution3D_CP_1129_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	226 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	368 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570__exit__
      -- CP-element group 232: 	 branch_block_stmt_453/getRemainingElementsx_xexit377_ifx_xend227
      -- CP-element group 232: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/$exit
      -- CP-element group 232: 	 branch_block_stmt_453/getRemainingElementsx_xexit377_ifx_xend227_PhiReq/$entry
      -- CP-element group 232: 	 branch_block_stmt_453/getRemainingElementsx_xexit377_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(226) & convolution3D_CP_1129_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	368 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Sample/cra
      -- 
    cra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1575_call_ack_0, ack => convolution3D_CP_1129_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	368 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	239 
    -- CP-element group 234: 	240 
    -- CP-element group 234: 	241 
    -- CP-element group 234: 	242 
    -- CP-element group 234: 	243 
    -- CP-element group 234: 	244 
    -- CP-element group 234:  members (28) 
      -- CP-element group 234: 	 branch_block_stmt_453/call_stmt_1575__exit__
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640__entry__
      -- CP-element group 234: 	 branch_block_stmt_453/call_stmt_1575/$exit
      -- CP-element group 234: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Update/cca
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_update_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_update_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_update_start_
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Update/cr
      -- 
    cca_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1575_call_ack_1, ack => convolution3D_CP_1129_elements(234)); -- 
    req_3078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => WPIPE_maxpool_output_pipe_1582_inst_req_0); -- 
    rr_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1615_inst_req_0); -- 
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1615_inst_req_1); -- 
    rr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1625_inst_req_0); -- 
    cr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1625_inst_req_1); -- 
    rr_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1634_inst_req_0); -- 
    cr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(234), ack => type_cast_1634_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_update_start_
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Update/req
      -- 
    ack_3079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_0, ack => convolution3D_CP_1129_elements(235)); -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(235), ack => WPIPE_maxpool_output_pipe_1582_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1582_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Sample/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_1, ack => convolution3D_CP_1129_elements(236)); -- 
    req_3092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(236), ack => WPIPE_maxpool_output_pipe_1586_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_update_start_
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Update/req
      -- 
    ack_3093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1586_inst_ack_0, ack => convolution3D_CP_1129_elements(237)); -- 
    req_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(237), ack => WPIPE_maxpool_output_pipe_1586_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	245 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/WPIPE_maxpool_output_pipe_1586_Update/ack
      -- 
    ack_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1586_inst_ack_1, ack => convolution3D_CP_1129_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	234 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Sample/ra
      -- 
    ra_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_0, ack => convolution3D_CP_1129_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	234 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	245 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1615_Update/ca
      -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_1, ack => convolution3D_CP_1129_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	234 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Sample/ra
      -- 
    ra_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => convolution3D_CP_1129_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	234 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	245 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1625_Update/ca
      -- 
    ca_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => convolution3D_CP_1129_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	234 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Sample/ra
      -- 
    ra_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_0, ack => convolution3D_CP_1129_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	234 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/type_cast_1634_Update/ca
      -- 
    ca_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_1, ack => convolution3D_CP_1129_elements(244)); -- 
    -- CP-element group 245:  join  transition  place  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	238 
    -- CP-element group 245: 	240 
    -- CP-element group 245: 	242 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	369 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640__exit__
      -- CP-element group 245: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody
      -- CP-element group 245: 	 branch_block_stmt_453/assign_stmt_1581_to_assign_stmt_1640/$exit
      -- CP-element group 245: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 245: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/$entry
      -- CP-element group 245: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/$entry
      -- 
    convolution3D_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(238) & convolution3D_CP_1129_elements(240) & convolution3D_CP_1129_elements(242) & convolution3D_CP_1129_elements(244);
      gj_convolution3D_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	374 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Sample/ra
      -- 
    ra_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_0, ack => convolution3D_CP_1129_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	374 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	254 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Update/ca
      -- 
    ca_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_1, ack => convolution3D_CP_1129_elements(247)); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	374 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_update_start_
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Sample/ack
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Update/req
      -- 
    ack_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1665_inst_ack_0, ack => convolution3D_CP_1129_elements(248)); -- 
    req_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(248), ack => WPIPE_num_out_pipe_1665_inst_req_1); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	259 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Update/ack
      -- 
    ack_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1665_inst_ack_1, ack => convolution3D_CP_1129_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	374 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Sample/ra
      -- 
    ra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_0, ack => convolution3D_CP_1129_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	374 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	254 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Update/ca
      -- 
    ca_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1670_inst_ack_1, ack => convolution3D_CP_1129_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	374 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Sample/ra
      -- 
    ra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_0, ack => convolution3D_CP_1129_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	374 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Update/ca
      -- 
    ca_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1674_inst_ack_1, ack => convolution3D_CP_1129_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	247 
    -- CP-element group 254: 	251 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Sample/crr
      -- 
    crr_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(254), ack => call_stmt_1685_call_req_0); -- 
    convolution3D_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(247) & convolution3D_CP_1129_elements(251) & convolution3D_CP_1129_elements(253);
      gj_convolution3D_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Sample/cra
      -- 
    cra_3208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_0, ack => convolution3D_CP_1129_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	374 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	259 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Update/cca
      -- 
    cca_3213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_1, ack => convolution3D_CP_1129_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	374 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Sample/cra
      -- 
    cra_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1692_call_ack_0, ack => convolution3D_CP_1129_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	374 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Update/cca
      -- 
    cca_3227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1692_call_ack_1, ack => convolution3D_CP_1129_elements(258)); -- 
    -- CP-element group 259:  branch  join  transition  place  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	249 
    -- CP-element group 259: 	256 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (10) 
      -- CP-element group 259: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703__exit__
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704__entry__
      -- CP-element group 259: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/$exit
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_dead_link/$entry
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_eval_test/$entry
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_eval_test/$exit
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_eval_test/branch_req
      -- CP-element group 259: 	 branch_block_stmt_453/R_exitcond5_1705_place
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_if_link/$entry
      -- CP-element group 259: 	 branch_block_stmt_453/if_stmt_1704_else_link/$entry
      -- 
    branch_req_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(259), ack => if_stmt_1704_branch_req_0); -- 
    convolution3D_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(249) & convolution3D_CP_1129_elements(256) & convolution3D_CP_1129_elements(258);
      gj_convolution3D_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: 	263 
    -- CP-element group 260:  members (18) 
      -- CP-element group 260: 	 branch_block_stmt_453/merge_stmt_1710__exit__
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715__entry__
      -- CP-element group 260: 	 branch_block_stmt_453/if_stmt_1704_if_link/$exit
      -- CP-element group 260: 	 branch_block_stmt_453/if_stmt_1704_if_link/if_choice_transition
      -- CP-element group 260: 	 branch_block_stmt_453/whilex_xbody_whilex_xend
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/$entry
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_update_start_
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_453/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 260: 	 branch_block_stmt_453/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 260: 	 branch_block_stmt_453/merge_stmt_1710_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_453/merge_stmt_1710_PhiAck/$entry
      -- CP-element group 260: 	 branch_block_stmt_453/merge_stmt_1710_PhiAck/$exit
      -- CP-element group 260: 	 branch_block_stmt_453/merge_stmt_1710_PhiAck/dummy
      -- 
    if_choice_transition_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1704_branch_ack_1, ack => convolution3D_CP_1129_elements(260)); -- 
    rr_3257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(260), ack => type_cast_1714_inst_req_0); -- 
    cr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(260), ack => type_cast_1714_inst_req_1); -- 
    -- CP-element group 261:  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	370 
    -- CP-element group 261: 	371 
    -- CP-element group 261:  members (12) 
      -- CP-element group 261: 	 branch_block_stmt_453/if_stmt_1704_else_link/$exit
      -- CP-element group 261: 	 branch_block_stmt_453/if_stmt_1704_else_link/else_choice_transition
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1704_branch_ack_0, ack => convolution3D_CP_1129_elements(261)); -- 
    rr_4028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(261), ack => type_cast_1646_inst_req_0); -- 
    cr_4033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(261), ack => type_cast_1646_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Sample/ra
      -- 
    ra_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1714_inst_ack_0, ack => convolution3D_CP_1129_elements(262)); -- 
    -- CP-element group 263:  fork  transition  place  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	260 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263: 	265 
    -- CP-element group 263: 	267 
    -- CP-element group 263: 	269 
    -- CP-element group 263: 	271 
    -- CP-element group 263: 	273 
    -- CP-element group 263: 	275 
    -- CP-element group 263: 	277 
    -- CP-element group 263: 	279 
    -- CP-element group 263: 	281 
    -- CP-element group 263: 	283 
    -- CP-element group 263:  members (40) 
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/assign_stmt_1715__exit__
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826__entry__
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/assign_stmt_1715/$exit
      -- CP-element group 263: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_453/assign_stmt_1715/type_cast_1714_Update/ca
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Sample/crr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Update/ccr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_update_start_
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Update/cr
      -- 
    ca_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1714_inst_ack_1, ack => convolution3D_CP_1129_elements(263)); -- 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1751_inst_req_1); -- 
    cr_3391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1791_inst_req_1); -- 
    cr_3349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1761_inst_req_1); -- 
    cr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1781_inst_req_1); -- 
    cr_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1801_inst_req_1); -- 
    cr_3363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1771_inst_req_1); -- 
    crr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => call_stmt_1718_call_req_0); -- 
    ccr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => call_stmt_1718_call_req_1); -- 
    cr_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1722_inst_req_1); -- 
    cr_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1731_inst_req_1); -- 
    cr_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(263), ack => type_cast_1741_inst_req_1); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Sample/cra
      -- 
    cra_3275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1718_call_ack_0, ack => convolution3D_CP_1129_elements(264)); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/call_stmt_1718_Update/cca
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Sample/rr
      -- 
    cca_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1718_call_ack_1, ack => convolution3D_CP_1129_elements(265)); -- 
    rr_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(265), ack => type_cast_1722_inst_req_0); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Sample/ra
      -- 
    ra_3289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1722_inst_ack_0, ack => convolution3D_CP_1129_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	263 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267: 	270 
    -- CP-element group 267: 	272 
    -- CP-element group 267: 	274 
    -- CP-element group 267: 	276 
    -- CP-element group 267: 	278 
    -- CP-element group 267: 	280 
    -- CP-element group 267: 	282 
    -- CP-element group 267:  members (27) 
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1722_Update/ca
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_sample_start_
      -- 
    ca_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1722_inst_ack_1, ack => convolution3D_CP_1129_elements(267)); -- 
    rr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1731_inst_req_0); -- 
    rr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1741_inst_req_0); -- 
    rr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1751_inst_req_0); -- 
    rr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1761_inst_req_0); -- 
    rr_3358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1771_inst_req_0); -- 
    rr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1781_inst_req_0); -- 
    rr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1791_inst_req_0); -- 
    rr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(267), ack => type_cast_1801_inst_req_0); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Sample/ra
      -- 
    ra_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_0, ack => convolution3D_CP_1129_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	263 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	304 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1731_Update/ca
      -- 
    ca_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_1, ack => convolution3D_CP_1129_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	267 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Sample/ra
      -- 
    ra_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_0, ack => convolution3D_CP_1129_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	263 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	301 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1741_Update/ca
      -- 
    ca_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1741_inst_ack_1, ack => convolution3D_CP_1129_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	267 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Sample/ra
      -- CP-element group 272: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_sample_completed_
      -- 
    ra_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1751_inst_ack_0, ack => convolution3D_CP_1129_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	263 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	298 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Update/ca
      -- CP-element group 273: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1751_update_completed_
      -- 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1751_inst_ack_1, ack => convolution3D_CP_1129_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	267 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Sample/$exit
      -- 
    ra_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1761_inst_ack_0, ack => convolution3D_CP_1129_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	263 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	295 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1761_update_completed_
      -- 
    ca_3350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1761_inst_ack_1, ack => convolution3D_CP_1129_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	267 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Sample/ra
      -- CP-element group 276: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_sample_completed_
      -- 
    ra_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1771_inst_ack_0, ack => convolution3D_CP_1129_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	263 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	292 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Update/ca
      -- CP-element group 277: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1771_Update/$exit
      -- 
    ca_3364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1771_inst_ack_1, ack => convolution3D_CP_1129_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	267 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Sample/ra
      -- CP-element group 278: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_sample_completed_
      -- 
    ra_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_0, ack => convolution3D_CP_1129_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	263 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	289 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Update/ca
      -- CP-element group 279: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1781_update_completed_
      -- 
    ca_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_1, ack => convolution3D_CP_1129_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	267 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Sample/ra
      -- CP-element group 280: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Sample/$exit
      -- 
    ra_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_0, ack => convolution3D_CP_1129_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	263 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	286 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Update/ca
      -- CP-element group 281: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1791_Update/$exit
      -- 
    ca_3392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_1, ack => convolution3D_CP_1129_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	267 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Sample/ra
      -- CP-element group 282: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_sample_completed_
      -- 
    ra_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_0, ack => convolution3D_CP_1129_elements(282)); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	263 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Update/ca
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/type_cast_1801_update_completed_
      -- 
    ca_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_1, ack => convolution3D_CP_1129_elements(283)); -- 
    req_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(283), ack => WPIPE_maxpool_output_pipe_1803_inst_req_0); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Update/req
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_update_start_
      -- CP-element group 284: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_sample_completed_
      -- 
    ack_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1803_inst_ack_0, ack => convolution3D_CP_1129_elements(284)); -- 
    req_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(284), ack => WPIPE_maxpool_output_pipe_1803_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1803_update_completed_
      -- 
    ack_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1803_inst_ack_1, ack => convolution3D_CP_1129_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	281 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_sample_start_
      -- 
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(286), ack => WPIPE_maxpool_output_pipe_1806_inst_req_0); -- 
    convolution3D_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(281) & convolution3D_CP_1129_elements(285);
      gj_convolution3D_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Update/req
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_update_start_
      -- CP-element group 287: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_sample_completed_
      -- 
    ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1806_inst_ack_0, ack => convolution3D_CP_1129_elements(287)); -- 
    req_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(287), ack => WPIPE_maxpool_output_pipe_1806_inst_req_1); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1806_update_completed_
      -- 
    ack_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1806_inst_ack_1, ack => convolution3D_CP_1129_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	279 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_sample_start_
      -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(289), ack => WPIPE_maxpool_output_pipe_1809_inst_req_0); -- 
    convolution3D_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(279) & convolution3D_CP_1129_elements(288);
      gj_convolution3D_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Update/req
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Sample/ack
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_update_start_
      -- CP-element group 290: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_sample_completed_
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1809_inst_ack_0, ack => convolution3D_CP_1129_elements(290)); -- 
    req_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(290), ack => WPIPE_maxpool_output_pipe_1809_inst_req_1); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Update/ack
      -- CP-element group 291: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1809_update_completed_
      -- 
    ack_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1809_inst_ack_1, ack => convolution3D_CP_1129_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	277 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Sample/req
      -- 
    req_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(292), ack => WPIPE_maxpool_output_pipe_1812_inst_req_0); -- 
    convolution3D_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(277) & convolution3D_CP_1129_elements(291);
      gj_convolution3D_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_update_start_
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Update/req
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Sample/$exit
      -- 
    ack_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1812_inst_ack_0, ack => convolution3D_CP_1129_elements(293)); -- 
    req_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(293), ack => WPIPE_maxpool_output_pipe_1812_inst_req_1); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1812_Update/$exit
      -- 
    ack_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1812_inst_ack_1, ack => convolution3D_CP_1129_elements(294)); -- 
    -- CP-element group 295:  join  transition  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	275 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_sample_start_
      -- 
    req_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(295), ack => WPIPE_maxpool_output_pipe_1815_inst_req_0); -- 
    convolution3D_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(275) & convolution3D_CP_1129_elements(294);
      gj_convolution3D_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Update/req
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Update/$entry
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Sample/ack
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_update_start_
      -- CP-element group 296: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_sample_completed_
      -- 
    ack_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1815_inst_ack_0, ack => convolution3D_CP_1129_elements(296)); -- 
    req_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(296), ack => WPIPE_maxpool_output_pipe_1815_inst_req_1); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1815_Update/ack
      -- 
    ack_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1815_inst_ack_1, ack => convolution3D_CP_1129_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	273 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_sample_start_
      -- 
    req_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(298), ack => WPIPE_maxpool_output_pipe_1818_inst_req_0); -- 
    convolution3D_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(273) & convolution3D_CP_1129_elements(297);
      gj_convolution3D_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Update/req
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_update_start_
      -- CP-element group 299: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_sample_completed_
      -- 
    ack_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1818_inst_ack_0, ack => convolution3D_CP_1129_elements(299)); -- 
    req_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(299), ack => WPIPE_maxpool_output_pipe_1818_inst_req_1); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1818_update_completed_
      -- 
    ack_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1818_inst_ack_1, ack => convolution3D_CP_1129_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	271 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_sample_start_
      -- 
    req_3498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(301), ack => WPIPE_maxpool_output_pipe_1821_inst_req_0); -- 
    convolution3D_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(271) & convolution3D_CP_1129_elements(300);
      gj_convolution3D_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Update/req
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Sample/ack
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Sample/$exit
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_update_start_
      -- CP-element group 302: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_sample_completed_
      -- 
    ack_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1821_inst_ack_0, ack => convolution3D_CP_1129_elements(302)); -- 
    req_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(302), ack => WPIPE_maxpool_output_pipe_1821_inst_req_1); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Update/ack
      -- CP-element group 303: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_Update/$exit
      -- CP-element group 303: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1821_update_completed_
      -- 
    ack_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1821_inst_ack_1, ack => convolution3D_CP_1129_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	269 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_sample_start_
      -- 
    req_3512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(304), ack => WPIPE_maxpool_output_pipe_1824_inst_req_0); -- 
    convolution3D_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(269) & convolution3D_CP_1129_elements(303);
      gj_convolution3D_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Update/req
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_update_start_
      -- CP-element group 305: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_sample_completed_
      -- 
    ack_3513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1824_inst_ack_0, ack => convolution3D_CP_1129_elements(305)); -- 
    req_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(305), ack => WPIPE_maxpool_output_pipe_1824_inst_req_1); -- 
    -- CP-element group 306:  transition  place  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (16) 
      -- CP-element group 306: 	 $exit
      -- CP-element group 306: 	 branch_block_stmt_453/$exit
      -- CP-element group 306: 	 branch_block_stmt_453/branch_block_stmt_453__exit__
      -- CP-element group 306: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826__exit__
      -- CP-element group 306: 	 branch_block_stmt_453/return__
      -- CP-element group 306: 	 branch_block_stmt_453/merge_stmt_1829__exit__
      -- CP-element group 306: 	 branch_block_stmt_453/merge_stmt_1829_PhiReqMerge
      -- CP-element group 306: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/WPIPE_maxpool_output_pipe_1824_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_453/call_stmt_1718_to_assign_stmt_1826/$exit
      -- CP-element group 306: 	 branch_block_stmt_453/return___PhiReq/$entry
      -- CP-element group 306: 	 branch_block_stmt_453/return___PhiReq/$exit
      -- CP-element group 306: 	 branch_block_stmt_453/merge_stmt_1829_PhiAck/$entry
      -- CP-element group 306: 	 branch_block_stmt_453/merge_stmt_1829_PhiAck/$exit
      -- CP-element group 306: 	 branch_block_stmt_453/merge_stmt_1829_PhiAck/dummy
      -- 
    ack_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1824_inst_ack_1, ack => convolution3D_CP_1129_elements(306)); -- 
    -- CP-element group 307:  transition  output  delay-element  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	86 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	311 
    -- CP-element group 307:  members (5) 
      -- CP-element group 307: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_req
      -- CP-element group 307: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_769_konst_delay_trans
      -- CP-element group 307: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/phi_stmt_763/$exit
      -- CP-element group 307: 	 branch_block_stmt_453/bbx_xnph389_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_763_req_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_763_req_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(307), ack => phi_stmt_763_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(307) is a control-delay.
    cp_element_307_delay: control_delay_element  generic map(name => " 307_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(86), ack => convolution3D_CP_1129_elements(307), clk => clk, reset =>reset);
    -- CP-element group 308:  transition  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	128 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Sample/ra
      -- CP-element group 308: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Sample/$exit
      -- 
    ra_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_0, ack => convolution3D_CP_1129_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	128 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (2) 
      -- CP-element group 309: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Update/ca
      -- CP-element group 309: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/Update/$exit
      -- 
    ca_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_1, ack => convolution3D_CP_1129_elements(309)); -- 
    -- CP-element group 310:  join  transition  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/SplitProtocol/$exit
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/type_cast_766/$exit
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_sources/$exit
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/$exit
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 310: 	 branch_block_stmt_453/forx_xbody_forx_xbody_PhiReq/phi_stmt_763/phi_stmt_763_req
      -- 
    phi_stmt_763_req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_763_req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(310), ack => phi_stmt_763_req_0); -- 
    convolution3D_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(308) & convolution3D_CP_1129_elements(309);
      gj_convolution3D_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  merge  transition  place  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	307 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (2) 
      -- CP-element group 311: 	 branch_block_stmt_453/merge_stmt_762_PhiAck/$entry
      -- CP-element group 311: 	 branch_block_stmt_453/merge_stmt_762_PhiReqMerge
      -- 
    convolution3D_CP_1129_elements(311) <= OrReduce(convolution3D_CP_1129_elements(307) & convolution3D_CP_1129_elements(310));
    -- CP-element group 312:  fork  transition  place  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	87 
    -- CP-element group 312: 	88 
    -- CP-element group 312: 	90 
    -- CP-element group 312: 	91 
    -- CP-element group 312: 	94 
    -- CP-element group 312: 	98 
    -- CP-element group 312: 	102 
    -- CP-element group 312: 	106 
    -- CP-element group 312: 	110 
    -- CP-element group 312: 	114 
    -- CP-element group 312: 	118 
    -- CP-element group 312: 	122 
    -- CP-element group 312: 	125 
    -- CP-element group 312:  members (56) 
      -- CP-element group 312: 	 branch_block_stmt_453/merge_stmt_762__exit__
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925__entry__
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_resized_1
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_scaled_1
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_computed_1
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_resize_1/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_resize_1/$exit
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_resize_1/index_resize_req
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_resize_1/index_resize_ack
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_scale_1/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_scale_1/$exit
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_scale_1/scale_rename_req
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_index_scale_1/scale_rename_ack
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_update_start
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Sample/req
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/array_obj_ref_775_final_index_sum_regn_Update/req
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_complete/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/addr_of_776_complete/req
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/RPIPE_maxpool_input_pipe_779_Sample/rr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_783_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_796_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_814_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_832_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_850_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_868_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_886_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/type_cast_904_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_update_start_
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/word_0/$entry
      -- CP-element group 312: 	 branch_block_stmt_453/assign_stmt_777_to_assign_stmt_925/ptr_deref_912_Update/word_access_complete/word_0/cr
      -- CP-element group 312: 	 branch_block_stmt_453/merge_stmt_762_PhiAck/phi_stmt_763_ack
      -- CP-element group 312: 	 branch_block_stmt_453/merge_stmt_762_PhiAck/$exit
      -- 
    phi_stmt_763_ack_3572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_763_ack_0, ack => convolution3D_CP_1129_elements(312)); -- 
    req_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => array_obj_ref_775_index_offset_req_0); -- 
    req_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => array_obj_ref_775_index_offset_req_1); -- 
    req_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => addr_of_776_final_reg_req_1); -- 
    rr_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => RPIPE_maxpool_input_pipe_779_inst_req_0); -- 
    cr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_783_inst_req_1); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_796_inst_req_1); -- 
    cr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_814_inst_req_1); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_832_inst_req_1); -- 
    cr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_850_inst_req_1); -- 
    cr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_868_inst_req_1); -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_886_inst_req_1); -- 
    cr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => type_cast_904_inst_req_1); -- 
    cr_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(312), ack => ptr_deref_912_store_0_req_1); -- 
    -- CP-element group 313:  transition  output  delay-element  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	76 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	317 
    -- CP-element group 313:  members (5) 
      -- CP-element group 313: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_req
      -- CP-element group 313: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_963_konst_delay_trans
      -- CP-element group 313: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/$exit
      -- CP-element group 313: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/phi_stmt_957/$exit
      -- CP-element group 313: 	 branch_block_stmt_453/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_957_req_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_957_req_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(313), ack => phi_stmt_957_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(313) is a control-delay.
    cp_element_313_delay: control_delay_element  generic map(name => " 313_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(76), ack => convolution3D_CP_1129_elements(313), clk => clk, reset =>reset);
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	127 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Sample/ra
      -- 
    ra_3615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_960_inst_ack_0, ack => convolution3D_CP_1129_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	127 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Update/ca
      -- CP-element group 315: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/Update/$exit
      -- 
    ca_3620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_960_inst_ack_1, ack => convolution3D_CP_1129_elements(315)); -- 
    -- CP-element group 316:  join  transition  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (6) 
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/SplitProtocol/$exit
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/type_cast_960/$exit
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_sources/$exit
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/$exit
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 316: 	 branch_block_stmt_453/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_957/phi_stmt_957_req
      -- 
    phi_stmt_957_req_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_957_req_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(316), ack => phi_stmt_957_req_0); -- 
    convolution3D_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(314) & convolution3D_CP_1129_elements(315);
      gj_convolution3D_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  merge  transition  place  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	313 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_453/merge_stmt_956_PhiReqMerge
      -- CP-element group 317: 	 branch_block_stmt_453/merge_stmt_956_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(317) <= OrReduce(convolution3D_CP_1129_elements(313) & convolution3D_CP_1129_elements(316));
    -- CP-element group 318:  branch  transition  place  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	129 
    -- CP-element group 318: 	130 
    -- CP-element group 318:  members (15) 
      -- CP-element group 318: 	 branch_block_stmt_453/merge_stmt_956__exit__
      -- CP-element group 318: 	 branch_block_stmt_453/assign_stmt_970_to_assign_stmt_976__entry__
      -- CP-element group 318: 	 branch_block_stmt_453/assign_stmt_970_to_assign_stmt_976__exit__
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977__entry__
      -- CP-element group 318: 	 branch_block_stmt_453/assign_stmt_970_to_assign_stmt_976/$entry
      -- CP-element group 318: 	 branch_block_stmt_453/assign_stmt_970_to_assign_stmt_976/$exit
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_dead_link/$entry
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_eval_test/$entry
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_eval_test/$exit
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_eval_test/branch_req
      -- CP-element group 318: 	 branch_block_stmt_453/R_tobool_978_place
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_if_link/$entry
      -- CP-element group 318: 	 branch_block_stmt_453/if_stmt_977_else_link/$entry
      -- CP-element group 318: 	 branch_block_stmt_453/merge_stmt_956_PhiAck/phi_stmt_957_ack
      -- CP-element group 318: 	 branch_block_stmt_453/merge_stmt_956_PhiAck/$exit
      -- 
    phi_stmt_957_ack_3626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_957_ack_0, ack => convolution3D_CP_1129_elements(318)); -- 
    branch_req_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(318), ack => if_stmt_977_branch_req_0); -- 
    -- CP-element group 319:  transition  output  delay-element  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	130 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (4) 
      -- CP-element group 319: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/$exit
      -- CP-element group 319: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1002_konst_delay_trans
      -- CP-element group 319: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_req
      -- CP-element group 319: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/$exit
      -- 
    phi_stmt_998_req_3649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_998_req_3649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(319), ack => phi_stmt_998_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(319) is a control-delay.
    cp_element_319_delay: control_delay_element  generic map(name => " 319_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(130), ack => convolution3D_CP_1129_elements(319), clk => clk, reset =>reset);
    -- CP-element group 320:  transition  output  delay-element  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	130 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (4) 
      -- CP-element group 320: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/$exit
      -- CP-element group 320: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/$exit
      -- CP-element group 320: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_req
      -- CP-element group 320: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1009_konst_delay_trans
      -- 
    phi_stmt_1005_req_3657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1005_req_3657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(320), ack => phi_stmt_1005_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(320) is a control-delay.
    cp_element_320_delay: control_delay_element  generic map(name => " 320_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(130), ack => convolution3D_CP_1129_elements(320), clk => clk, reset =>reset);
    -- CP-element group 321:  join  transition  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	329 
    -- CP-element group 321:  members (1) 
      -- CP-element group 321: 	 branch_block_stmt_453/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(319) & convolution3D_CP_1129_elements(320);
      gj_convolution3D_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	138 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Sample/ra
      -- 
    ra_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_0, ack => convolution3D_CP_1129_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	138 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Update/ca
      -- CP-element group 323: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/Update/$exit
      -- 
    ca_3682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_1, ack => convolution3D_CP_1129_elements(323)); -- 
    -- CP-element group 324:  join  transition  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	328 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/SplitProtocol/$exit
      -- CP-element group 324: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/type_cast_1004/$exit
      -- CP-element group 324: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_req
      -- CP-element group 324: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/phi_stmt_998_sources/$exit
      -- CP-element group 324: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_998/$exit
      -- 
    phi_stmt_998_req_3683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_998_req_3683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(324), ack => phi_stmt_998_req_1); -- 
    convolution3D_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(322) & convolution3D_CP_1129_elements(323);
      gj_convolution3D_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	138 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (2) 
      -- CP-element group 325: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Sample/ra
      -- CP-element group 325: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Sample/$exit
      -- 
    ra_3700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1011_inst_ack_0, ack => convolution3D_CP_1129_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	138 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (2) 
      -- CP-element group 326: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/Update/ca
      -- 
    ca_3705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1011_inst_ack_1, ack => convolution3D_CP_1129_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/SplitProtocol/$exit
      -- CP-element group 327: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/type_cast_1011/$exit
      -- CP-element group 327: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/$exit
      -- CP-element group 327: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1005/phi_stmt_1005_req
      -- 
    phi_stmt_1005_req_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1005_req_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(327), ack => phi_stmt_1005_req_1); -- 
    convolution3D_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(325) & convolution3D_CP_1129_elements(326);
      gj_convolution3D_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	324 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_453/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(324) & convolution3D_CP_1129_elements(327);
      gj_convolution3D_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  merge  fork  transition  place  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	321 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_453/merge_stmt_997_PhiReqMerge
      -- CP-element group 329: 	 branch_block_stmt_453/merge_stmt_997_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(329) <= OrReduce(convolution3D_CP_1129_elements(321) & convolution3D_CP_1129_elements(328));
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_453/merge_stmt_997_PhiAck/phi_stmt_998_ack
      -- 
    phi_stmt_998_ack_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_998_ack_0, ack => convolution3D_CP_1129_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (1) 
      -- CP-element group 331: 	 branch_block_stmt_453/merge_stmt_997_PhiAck/phi_stmt_1005_ack
      -- 
    phi_stmt_1005_ack_3712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1005_ack_0, ack => convolution3D_CP_1129_elements(331)); -- 
    -- CP-element group 332:  join  fork  transition  place  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	131 
    -- CP-element group 332: 	134 
    -- CP-element group 332: 	135 
    -- CP-element group 332: 	136 
    -- CP-element group 332:  members (16) 
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_update_start_
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Sample/rr
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Update/$entry
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_Update/cr
      -- CP-element group 332: 	 branch_block_stmt_453/merge_stmt_997__exit__
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051__entry__
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1045_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/$entry
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/RPIPE_maxpool_input_pipe_1026_Sample/rr
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_update_start_
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Update/$entry
      -- CP-element group 332: 	 branch_block_stmt_453/assign_stmt_1018_to_assign_stmt_1051/type_cast_1030_Update/cr
      -- CP-element group 332: 	 branch_block_stmt_453/merge_stmt_997_PhiAck/$exit
      -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(332), ack => type_cast_1045_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(332), ack => type_cast_1045_inst_req_1); -- 
    rr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(332), ack => RPIPE_maxpool_input_pipe_1026_inst_req_0); -- 
    cr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(332), ack => type_cast_1030_inst_req_1); -- 
    convolution3D_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(330) & convolution3D_CP_1129_elements(331);
      gj_convolution3D_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	139 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Sample/ra
      -- 
    ra_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_0, ack => convolution3D_CP_1129_elements(333)); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	139 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/Update/ca
      -- 
    ca_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1062_inst_ack_1, ack => convolution3D_CP_1129_elements(334)); -- 
    -- CP-element group 335:  join  transition  place  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (8) 
      -- CP-element group 335: 	 branch_block_stmt_453/merge_stmt_1058_PhiReqMerge
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/$exit
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$exit
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/$exit
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1062/SplitProtocol/$exit
      -- CP-element group 335: 	 branch_block_stmt_453/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1059/phi_stmt_1059_req
      -- CP-element group 335: 	 branch_block_stmt_453/merge_stmt_1058_PhiAck/$entry
      -- 
    phi_stmt_1059_req_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_req_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(335), ack => phi_stmt_1059_req_0); -- 
    convolution3D_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(333) & convolution3D_CP_1129_elements(334);
      gj_convolution3D_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	140 
    -- CP-element group 336: 	141 
    -- CP-element group 336: 	143 
    -- CP-element group 336: 	145 
    -- CP-element group 336:  members (29) 
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_update_start_
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Update/req
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Update/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_complete/req
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/word_0/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_Update/word_access_complete/word_0/cr
      -- CP-element group 336: 	 branch_block_stmt_453/merge_stmt_1058__exit__
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097__entry__
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_resized_1
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_scaled_1
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_computed_1
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Sample/req
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_final_index_sum_regn_update_start
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_scale_1/scale_rename_ack
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_scale_1/scale_rename_req
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_scale_1/$exit
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_scale_1/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_resize_1/index_resize_ack
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_resize_1/index_resize_req
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_resize_1/$exit
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/addr_of_1092_complete/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/ptr_deref_1095_update_start_
      -- CP-element group 336: 	 branch_block_stmt_453/assign_stmt_1069_to_assign_stmt_1097/array_obj_ref_1091_index_resize_1/$entry
      -- CP-element group 336: 	 branch_block_stmt_453/merge_stmt_1058_PhiAck/$exit
      -- CP-element group 336: 	 branch_block_stmt_453/merge_stmt_1058_PhiAck/phi_stmt_1059_ack
      -- 
    phi_stmt_1059_ack_3747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1059_ack_0, ack => convolution3D_CP_1129_elements(336)); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(336), ack => array_obj_ref_1091_index_offset_req_1); -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(336), ack => addr_of_1092_final_reg_req_1); -- 
    cr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(336), ack => ptr_deref_1095_store_0_req_1); -- 
    req_2267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(336), ack => array_obj_ref_1091_index_offset_req_0); -- 
    -- CP-element group 337:  merge  fork  transition  place  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	129 
    -- CP-element group 337: 	146 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	147 
    -- CP-element group 337: 	148 
    -- CP-element group 337: 	149 
    -- CP-element group 337: 	150 
    -- CP-element group 337: 	151 
    -- CP-element group 337: 	152 
    -- CP-element group 337: 	153 
    -- CP-element group 337: 	154 
    -- CP-element group 337:  members (31) 
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_update_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_453/merge_stmt_1099_PhiReqMerge
      -- CP-element group 337: 	 branch_block_stmt_453/merge_stmt_1099__exit__
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151__entry__
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_update_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1114_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_update_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1110_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_update_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1102_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Sample/rr
      -- CP-element group 337: 	 branch_block_stmt_453/assign_stmt_1103_to_assign_stmt_1151/type_cast_1106_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/merge_stmt_1099_PhiAck/$entry
      -- CP-element group 337: 	 branch_block_stmt_453/merge_stmt_1099_PhiAck/$exit
      -- CP-element group 337: 	 branch_block_stmt_453/merge_stmt_1099_PhiAck/dummy
      -- 
    cr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1102_inst_req_1); -- 
    rr_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1102_inst_req_0); -- 
    cr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1114_inst_req_1); -- 
    rr_2391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1114_inst_req_0); -- 
    cr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1110_inst_req_1); -- 
    rr_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1110_inst_req_0); -- 
    cr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1106_inst_req_1); -- 
    rr_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(337), ack => type_cast_1106_inst_req_0); -- 
    convolution3D_CP_1129_elements(337) <= OrReduce(convolution3D_CP_1129_elements(129) & convolution3D_CP_1129_elements(146));
    -- CP-element group 338:  transition  output  delay-element  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	170 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	342 
    -- CP-element group 338:  members (5) 
      -- CP-element group 338: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 338: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/$exit
      -- CP-element group 338: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/$exit
      -- CP-element group 338: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1236_konst_delay_trans
      -- CP-element group 338: 	 branch_block_stmt_453/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_req
      -- 
    phi_stmt_1232_req_3781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1232_req_3781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(338), ack => phi_stmt_1232_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(338) is a control-delay.
    cp_element_338_delay: control_delay_element  generic map(name => " 338_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(170), ack => convolution3D_CP_1129_elements(338), clk => clk, reset =>reset);
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	212 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (2) 
      -- CP-element group 339: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Sample/ra
      -- 
    ra_3801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convolution3D_CP_1129_elements(339)); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	212 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/Update/ca
      -- 
    ca_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convolution3D_CP_1129_elements(340)); -- 
    -- CP-element group 341:  join  transition  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/$exit
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/$exit
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/$exit
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_sources/type_cast_1238/SplitProtocol/$exit
      -- CP-element group 341: 	 branch_block_stmt_453/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1232/phi_stmt_1232_req
      -- 
    phi_stmt_1232_req_3807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1232_req_3807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(341), ack => phi_stmt_1232_req_1); -- 
    convolution3D_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(339) & convolution3D_CP_1129_elements(340);
      gj_convolution3D_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  merge  transition  place  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	338 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (2) 
      -- CP-element group 342: 	 branch_block_stmt_453/merge_stmt_1231_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_453/merge_stmt_1231_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(342) <= OrReduce(convolution3D_CP_1129_elements(338) & convolution3D_CP_1129_elements(341));
    -- CP-element group 343:  fork  transition  place  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	171 
    -- CP-element group 343: 	172 
    -- CP-element group 343: 	174 
    -- CP-element group 343: 	175 
    -- CP-element group 343: 	178 
    -- CP-element group 343: 	182 
    -- CP-element group 343: 	186 
    -- CP-element group 343: 	190 
    -- CP-element group 343: 	194 
    -- CP-element group 343: 	198 
    -- CP-element group 343: 	202 
    -- CP-element group 343: 	206 
    -- CP-element group 343: 	209 
    -- CP-element group 343:  members (56) 
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_update_start
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Sample/req
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/merge_stmt_1231__exit__
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394__entry__
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_final_index_sum_regn_Update/req
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_scale_1/scale_rename_ack
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_scale_1/scale_rename_req
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_scale_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_scale_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_resize_1/index_resize_ack
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_resize_1/index_resize_req
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_resize_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_resize_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_computed_1
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_scaled_1
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1301_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/array_obj_ref_1244_index_resized_1
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1252_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1283_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Sample/rr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/RPIPE_maxpool_input_pipe_1248_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1265_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1319_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/addr_of_1245_complete/req
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1337_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1355_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/type_cast_1373_Update/cr
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_update_start_
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 branch_block_stmt_453/assign_stmt_1246_to_assign_stmt_1394/ptr_deref_1381_Update/word_access_complete/word_0/cr
      -- CP-element group 343: 	 branch_block_stmt_453/merge_stmt_1231_PhiAck/$exit
      -- CP-element group 343: 	 branch_block_stmt_453/merge_stmt_1231_PhiAck/phi_stmt_1232_ack
      -- 
    phi_stmt_1232_ack_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1232_ack_0, ack => convolution3D_CP_1129_elements(343)); -- 
    req_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => array_obj_ref_1244_index_offset_req_0); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => array_obj_ref_1244_index_offset_req_1); -- 
    cr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1301_inst_req_1); -- 
    cr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1252_inst_req_1); -- 
    cr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1265_inst_req_1); -- 
    cr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1283_inst_req_1); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1319_inst_req_1); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => RPIPE_maxpool_input_pipe_1248_inst_req_0); -- 
    req_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => addr_of_1245_final_reg_req_1); -- 
    cr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1337_inst_req_1); -- 
    cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1355_inst_req_1); -- 
    cr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => type_cast_1373_inst_req_1); -- 
    cr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(343), ack => ptr_deref_1381_store_0_req_1); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	211 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (2) 
      -- CP-element group 344: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Sample/ra
      -- 
    ra_3844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => convolution3D_CP_1129_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	211 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (2) 
      -- CP-element group 345: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/Update/ca
      -- 
    ca_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => convolution3D_CP_1129_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/$exit
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$exit
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/$exit
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1429/SplitProtocol/$exit
      -- CP-element group 346: 	 branch_block_stmt_453/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_req
      -- 
    phi_stmt_1426_req_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1426_req_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(346), ack => phi_stmt_1426_req_0); -- 
    convolution3D_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(344) & convolution3D_CP_1129_elements(345);
      gj_convolution3D_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  transition  output  delay-element  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	157 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (5) 
      -- CP-element group 347: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 347: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/$exit
      -- CP-element group 347: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$exit
      -- CP-element group 347: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432_konst_delay_trans
      -- CP-element group 347: 	 branch_block_stmt_453/ifx_xend_forx_xend215_PhiReq/phi_stmt_1426/phi_stmt_1426_req
      -- 
    phi_stmt_1426_req_3861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1426_req_3861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(347), ack => phi_stmt_1426_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(347) is a control-delay.
    cp_element_347_delay: control_delay_element  generic map(name => " 347_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(157), ack => convolution3D_CP_1129_elements(347), clk => clk, reset =>reset);
    -- CP-element group 348:  merge  transition  place  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (2) 
      -- CP-element group 348: 	 branch_block_stmt_453/merge_stmt_1425_PhiReqMerge
      -- CP-element group 348: 	 branch_block_stmt_453/merge_stmt_1425_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(348) <= OrReduce(convolution3D_CP_1129_elements(346) & convolution3D_CP_1129_elements(347));
    -- CP-element group 349:  branch  transition  place  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	213 
    -- CP-element group 349: 	214 
    -- CP-element group 349:  members (15) 
      -- CP-element group 349: 	 branch_block_stmt_453/merge_stmt_1425__exit__
      -- CP-element group 349: 	 branch_block_stmt_453/assign_stmt_1439_to_assign_stmt_1445__entry__
      -- CP-element group 349: 	 branch_block_stmt_453/assign_stmt_1439_to_assign_stmt_1445__exit__
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446__entry__
      -- CP-element group 349: 	 branch_block_stmt_453/assign_stmt_1439_to_assign_stmt_1445/$entry
      -- CP-element group 349: 	 branch_block_stmt_453/assign_stmt_1439_to_assign_stmt_1445/$exit
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_dead_link/$entry
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_eval_test/$entry
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_eval_test/$exit
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_eval_test/branch_req
      -- CP-element group 349: 	 branch_block_stmt_453/R_tobool218_1447_place
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_if_link/$entry
      -- CP-element group 349: 	 branch_block_stmt_453/if_stmt_1446_else_link/$entry
      -- CP-element group 349: 	 branch_block_stmt_453/merge_stmt_1425_PhiAck/$exit
      -- CP-element group 349: 	 branch_block_stmt_453/merge_stmt_1425_PhiAck/phi_stmt_1426_ack
      -- 
    phi_stmt_1426_ack_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1426_ack_0, ack => convolution3D_CP_1129_elements(349)); -- 
    branch_req_2859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(349), ack => if_stmt_1446_branch_req_0); -- 
    -- CP-element group 350:  transition  output  delay-element  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	216 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (4) 
      -- CP-element group 350: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/$exit
      -- CP-element group 350: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$exit
      -- CP-element group 350: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1475_konst_delay_trans
      -- CP-element group 350: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_req
      -- 
    phi_stmt_1471_req_3889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1471_req_3889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(350), ack => phi_stmt_1471_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(350) is a control-delay.
    cp_element_350_delay: control_delay_element  generic map(name => " 350_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(216), ack => convolution3D_CP_1129_elements(350), clk => clk, reset =>reset);
    -- CP-element group 351:  transition  output  delay-element  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	216 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (4) 
      -- CP-element group 351: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/$exit
      -- CP-element group 351: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/$exit
      -- CP-element group 351: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1482_konst_delay_trans
      -- CP-element group 351: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_req
      -- 
    phi_stmt_1478_req_3897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1478_req_3897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(351), ack => phi_stmt_1478_req_0); -- 
    -- Element group convolution3D_CP_1129_elements(351) is a control-delay.
    cp_element_351_delay: control_delay_element  generic map(name => " 351_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(216), ack => convolution3D_CP_1129_elements(351), clk => clk, reset =>reset);
    -- CP-element group 352:  join  transition  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	360 
    -- CP-element group 352:  members (1) 
      -- CP-element group 352: 	 branch_block_stmt_453/bbx_xnphx_xi360_forx_xbodyx_xi369_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(350) & convolution3D_CP_1129_elements(351);
      gj_convolution3D_cp_element_group_352 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	224 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (2) 
      -- CP-element group 353: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Sample/ra
      -- 
    ra_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1477_inst_ack_0, ack => convolution3D_CP_1129_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	224 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (2) 
      -- CP-element group 354: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/Update/ca
      -- 
    ca_3922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1477_inst_ack_1, ack => convolution3D_CP_1129_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	359 
    -- CP-element group 355:  members (5) 
      -- CP-element group 355: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/$exit
      -- CP-element group 355: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/$exit
      -- CP-element group 355: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/$exit
      -- CP-element group 355: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_sources/type_cast_1477/SplitProtocol/$exit
      -- CP-element group 355: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1471/phi_stmt_1471_req
      -- 
    phi_stmt_1471_req_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1471_req_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(355), ack => phi_stmt_1471_req_1); -- 
    convolution3D_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(353) & convolution3D_CP_1129_elements(354);
      gj_convolution3D_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	224 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (2) 
      -- CP-element group 356: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Sample/ra
      -- 
    ra_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1484_inst_ack_0, ack => convolution3D_CP_1129_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	224 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (2) 
      -- CP-element group 357: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/Update/ca
      -- 
    ca_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1484_inst_ack_1, ack => convolution3D_CP_1129_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (5) 
      -- CP-element group 358: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/$exit
      -- CP-element group 358: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/$exit
      -- CP-element group 358: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/$exit
      -- CP-element group 358: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_sources/type_cast_1484/SplitProtocol/$exit
      -- CP-element group 358: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/phi_stmt_1478/phi_stmt_1478_req
      -- 
    phi_stmt_1478_req_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1478_req_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(358), ack => phi_stmt_1478_req_1); -- 
    convolution3D_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(356) & convolution3D_CP_1129_elements(357);
      gj_convolution3D_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  join  transition  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	355 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (1) 
      -- CP-element group 359: 	 branch_block_stmt_453/forx_xbodyx_xi369_forx_xbodyx_xi369_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(355) & convolution3D_CP_1129_elements(358);
      gj_convolution3D_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  merge  fork  transition  place  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	352 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_453/merge_stmt_1470_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_453/merge_stmt_1470_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(360) <= OrReduce(convolution3D_CP_1129_elements(352) & convolution3D_CP_1129_elements(359));
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (1) 
      -- CP-element group 361: 	 branch_block_stmt_453/merge_stmt_1470_PhiAck/phi_stmt_1471_ack
      -- 
    phi_stmt_1471_ack_3951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1471_ack_0, ack => convolution3D_CP_1129_elements(361)); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (1) 
      -- CP-element group 362: 	 branch_block_stmt_453/merge_stmt_1470_PhiAck/phi_stmt_1478_ack
      -- 
    phi_stmt_1478_ack_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1478_ack_0, ack => convolution3D_CP_1129_elements(362)); -- 
    -- CP-element group 363:  join  fork  transition  place  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	217 
    -- CP-element group 363: 	220 
    -- CP-element group 363: 	221 
    -- CP-element group 363: 	222 
    -- CP-element group 363:  members (16) 
      -- CP-element group 363: 	 branch_block_stmt_453/merge_stmt_1470__exit__
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524__entry__
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/$entry
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/RPIPE_maxpool_input_pipe_1499_Sample/rr
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_update_start_
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1503_Update/cr
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_update_start_
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Sample/rr
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_453/assign_stmt_1491_to_assign_stmt_1524/type_cast_1518_Update/cr
      -- CP-element group 363: 	 branch_block_stmt_453/merge_stmt_1470_PhiAck/$exit
      -- 
    rr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(363), ack => RPIPE_maxpool_input_pipe_1499_inst_req_0); -- 
    cr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(363), ack => type_cast_1503_inst_req_1); -- 
    rr_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(363), ack => type_cast_1518_inst_req_0); -- 
    cr_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(363), ack => type_cast_1518_inst_req_1); -- 
    convolution3D_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(361) & convolution3D_CP_1129_elements(362);
      gj_convolution3D_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	225 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	366 
    -- CP-element group 364:  members (2) 
      -- CP-element group 364: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Sample/ra
      -- 
    ra_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_0, ack => convolution3D_CP_1129_elements(364)); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	225 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/Update/ca
      -- 
    ca_3981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_1, ack => convolution3D_CP_1129_elements(365)); -- 
    -- CP-element group 366:  join  transition  place  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	364 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (8) 
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/$exit
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/$exit
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/$exit
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/$exit
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_sources/type_cast_1535/SplitProtocol/$exit
      -- CP-element group 366: 	 branch_block_stmt_453/forx_xbodyx_xi369_getRemainingElementsx_xexit377_PhiReq/phi_stmt_1532/phi_stmt_1532_req
      -- CP-element group 366: 	 branch_block_stmt_453/merge_stmt_1531_PhiReqMerge
      -- CP-element group 366: 	 branch_block_stmt_453/merge_stmt_1531_PhiAck/$entry
      -- 
    phi_stmt_1532_req_3982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1532_req_3982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(366), ack => phi_stmt_1532_req_0); -- 
    convolution3D_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(364) & convolution3D_CP_1129_elements(365);
      gj_convolution3D_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	226 
    -- CP-element group 367: 	227 
    -- CP-element group 367: 	229 
    -- CP-element group 367: 	231 
    -- CP-element group 367:  members (29) 
      -- CP-element group 367: 	 branch_block_stmt_453/merge_stmt_1531__exit__
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570__entry__
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_update_start_
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_resized_1
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_scaled_1
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_computed_1
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_resize_1/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_resize_1/$exit
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_resize_1/index_resize_req
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_resize_1/index_resize_ack
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_scale_1/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_scale_1/$exit
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_scale_1/scale_rename_req
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_index_scale_1/scale_rename_ack
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_update_start
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Sample/req
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/array_obj_ref_1564_final_index_sum_regn_Update/req
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_complete/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/addr_of_1565_complete/req
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_update_start_
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/word_0/$entry
      -- CP-element group 367: 	 branch_block_stmt_453/assign_stmt_1542_to_assign_stmt_1570/ptr_deref_1568_Update/word_access_complete/word_0/cr
      -- CP-element group 367: 	 branch_block_stmt_453/merge_stmt_1531_PhiAck/$exit
      -- CP-element group 367: 	 branch_block_stmt_453/merge_stmt_1531_PhiAck/phi_stmt_1532_ack
      -- 
    phi_stmt_1532_ack_3987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1532_ack_0, ack => convolution3D_CP_1129_elements(367)); -- 
    req_2979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(367), ack => array_obj_ref_1564_index_offset_req_0); -- 
    req_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(367), ack => array_obj_ref_1564_index_offset_req_1); -- 
    req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(367), ack => addr_of_1565_final_reg_req_1); -- 
    cr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(367), ack => ptr_deref_1568_store_0_req_1); -- 
    -- CP-element group 368:  merge  fork  transition  place  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	213 
    -- CP-element group 368: 	232 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	233 
    -- CP-element group 368: 	234 
    -- CP-element group 368:  members (13) 
      -- CP-element group 368: 	 branch_block_stmt_453/merge_stmt_1572__exit__
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575__entry__
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/$entry
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_update_start_
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Sample/crr
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_453/call_stmt_1575/call_stmt_1575_Update/ccr
      -- CP-element group 368: 	 branch_block_stmt_453/merge_stmt_1572_PhiReqMerge
      -- CP-element group 368: 	 branch_block_stmt_453/merge_stmt_1572_PhiAck/$entry
      -- CP-element group 368: 	 branch_block_stmt_453/merge_stmt_1572_PhiAck/$exit
      -- CP-element group 368: 	 branch_block_stmt_453/merge_stmt_1572_PhiAck/dummy
      -- 
    crr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(368), ack => call_stmt_1575_call_req_0); -- 
    ccr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(368), ack => call_stmt_1575_call_req_1); -- 
    convolution3D_CP_1129_elements(368) <= OrReduce(convolution3D_CP_1129_elements(213) & convolution3D_CP_1129_elements(232));
    -- CP-element group 369:  transition  output  delay-element  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	245 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	373 
    -- CP-element group 369:  members (5) 
      -- CP-element group 369: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 369: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/$exit
      -- CP-element group 369: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/$exit
      -- CP-element group 369: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1649_konst_delay_trans
      -- CP-element group 369: 	 branch_block_stmt_453/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_req
      -- 
    phi_stmt_1643_req_4009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1643_req_4009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(369), ack => phi_stmt_1643_req_1); -- 
    -- Element group convolution3D_CP_1129_elements(369) is a control-delay.
    cp_element_369_delay: control_delay_element  generic map(name => " 369_delay", delay_value => 1)  port map(req => convolution3D_CP_1129_elements(245), ack => convolution3D_CP_1129_elements(369), clk => clk, reset =>reset);
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	261 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Sample/ra
      -- 
    ra_4029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_0, ack => convolution3D_CP_1129_elements(370)); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	261 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/Update/ca
      -- 
    ca_4034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_1, ack => convolution3D_CP_1129_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/$exit
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/$exit
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/$exit
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_sources/type_cast_1646/SplitProtocol/$exit
      -- CP-element group 372: 	 branch_block_stmt_453/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1643/phi_stmt_1643_req
      -- 
    phi_stmt_1643_req_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1643_req_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(372), ack => phi_stmt_1643_req_0); -- 
    convolution3D_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1129_elements(370) & convolution3D_CP_1129_elements(371);
      gj_convolution3D_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1129_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  merge  transition  place  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	369 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (2) 
      -- CP-element group 373: 	 branch_block_stmt_453/merge_stmt_1642_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_453/merge_stmt_1642_PhiAck/$entry
      -- 
    convolution3D_CP_1129_elements(373) <= OrReduce(convolution3D_CP_1129_elements(369) & convolution3D_CP_1129_elements(372));
    -- CP-element group 374:  fork  transition  place  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	246 
    -- CP-element group 374: 	247 
    -- CP-element group 374: 	248 
    -- CP-element group 374: 	250 
    -- CP-element group 374: 	251 
    -- CP-element group 374: 	252 
    -- CP-element group 374: 	253 
    -- CP-element group 374: 	256 
    -- CP-element group 374: 	257 
    -- CP-element group 374: 	258 
    -- CP-element group 374:  members (35) 
      -- CP-element group 374: 	 branch_block_stmt_453/merge_stmt_1642__exit__
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703__entry__
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_update_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Sample/rr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1663_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/WPIPE_num_out_pipe_1665_Sample/req
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_update_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Sample/rr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1670_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_update_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Sample/rr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/type_cast_1674_Update/cr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_update_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1685_Update/ccr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_update_start_
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Sample/crr
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_453/assign_stmt_1655_to_assign_stmt_1703/call_stmt_1692_Update/ccr
      -- CP-element group 374: 	 branch_block_stmt_453/merge_stmt_1642_PhiAck/$exit
      -- CP-element group 374: 	 branch_block_stmt_453/merge_stmt_1642_PhiAck/phi_stmt_1643_ack
      -- 
    phi_stmt_1643_ack_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1643_ack_0, ack => convolution3D_CP_1129_elements(374)); -- 
    rr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1663_inst_req_0); -- 
    cr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1663_inst_req_1); -- 
    req_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => WPIPE_num_out_pipe_1665_inst_req_0); -- 
    rr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1670_inst_req_0); -- 
    cr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1670_inst_req_1); -- 
    rr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1674_inst_req_0); -- 
    cr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => type_cast_1674_inst_req_1); -- 
    ccr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => call_stmt_1685_call_req_1); -- 
    crr_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => call_stmt_1692_call_req_0); -- 
    ccr_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1129_elements(374), ack => call_stmt_1692_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1143_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1421_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_952_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1069 : std_logic_vector(63 downto 0);
    signal R_indvar417_1243_resized : std_logic_vector(13 downto 0);
    signal R_indvar417_1243_scaled : std_logic_vector(13 downto 0);
    signal R_indvar431_774_resized : std_logic_vector(13 downto 0);
    signal R_indvar431_774_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1090_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1090_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1563_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1563_scaled : std_logic_vector(13 downto 0);
    signal add102_820 : std_logic_vector(63 downto 0);
    signal add108_838 : std_logic_vector(63 downto 0);
    signal add114_856 : std_logic_vector(63 downto 0);
    signal add120_874 : std_logic_vector(63 downto 0);
    signal add1216x_xi374_1548 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1075 : std_logic_vector(63 downto 0);
    signal add126_892 : std_logic_vector(63 downto 0);
    signal add132_910 : std_logic_vector(63 downto 0);
    signal add13_504 : std_logic_vector(15 downto 0);
    signal add171_1271 : std_logic_vector(63 downto 0);
    signal add177_1289 : std_logic_vector(63 downto 0);
    signal add183_1307 : std_logic_vector(63 downto 0);
    signal add189_1325 : std_logic_vector(63 downto 0);
    signal add195_1343 : std_logic_vector(63 downto 0);
    signal add201_1361 : std_logic_vector(63 downto 0);
    signal add207_1379 : std_logic_vector(63 downto 0);
    signal add23_529 : std_logic_vector(15 downto 0);
    signal add33_554 : std_logic_vector(15 downto 0);
    signal add43_579 : std_logic_vector(15 downto 0);
    signal add53_604 : std_logic_vector(15 downto 0);
    signal add63_629 : std_logic_vector(15 downto 0);
    signal add73_654 : std_logic_vector(15 downto 0);
    signal add96_802 : std_logic_vector(63 downto 0);
    signal add_479 : std_logic_vector(31 downto 0);
    signal addx_xi365_1509 : std_logic_vector(63 downto 0);
    signal addx_xi_1036 : std_logic_vector(63 downto 0);
    signal and217_1439 : std_logic_vector(63 downto 0);
    signal and264_1681 : std_logic_vector(7 downto 0);
    signal and_970 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1091_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1091_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1091_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1091_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1091_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1091_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1244_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1564_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_775_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1093 : std_logic_vector(31 downto 0);
    signal arrayidx211_1246 : std_logic_vector(31 downto 0);
    signal arrayidx226_1566 : std_logic_vector(31 downto 0);
    signal arrayidx_777 : std_logic_vector(31 downto 0);
    signal call105_829 : std_logic_vector(7 downto 0);
    signal call111_847 : std_logic_vector(7 downto 0);
    signal call117_865 : std_logic_vector(7 downto 0);
    signal call11_495 : std_logic_vector(7 downto 0);
    signal call123_883 : std_logic_vector(7 downto 0);
    signal call129_901 : std_logic_vector(7 downto 0);
    signal call164_1249 : std_logic_vector(7 downto 0);
    signal call168_1262 : std_logic_vector(7 downto 0);
    signal call16_507 : std_logic_vector(7 downto 0);
    signal call174_1280 : std_logic_vector(7 downto 0);
    signal call180_1298 : std_logic_vector(7 downto 0);
    signal call186_1316 : std_logic_vector(7 downto 0);
    signal call192_1334 : std_logic_vector(7 downto 0);
    signal call198_1352 : std_logic_vector(7 downto 0);
    signal call204_1370 : std_logic_vector(7 downto 0);
    signal call21_520 : std_logic_vector(7 downto 0);
    signal call229_1575 : std_logic_vector(63 downto 0);
    signal call26_532 : std_logic_vector(7 downto 0);
    signal call288_1718 : std_logic_vector(63 downto 0);
    signal call2_470 : std_logic_vector(7 downto 0);
    signal call31_545 : std_logic_vector(7 downto 0);
    signal call36_557 : std_logic_vector(7 downto 0);
    signal call41_570 : std_logic_vector(7 downto 0);
    signal call46_582 : std_logic_vector(7 downto 0);
    signal call51_595 : std_logic_vector(7 downto 0);
    signal call56_607 : std_logic_vector(7 downto 0);
    signal call61_620 : std_logic_vector(7 downto 0);
    signal call66_632 : std_logic_vector(7 downto 0);
    signal call6_482 : std_logic_vector(7 downto 0);
    signal call71_645 : std_logic_vector(7 downto 0);
    signal call89_780 : std_logic_vector(7 downto 0);
    signal call93_793 : std_logic_vector(7 downto 0);
    signal call99_811 : std_logic_vector(7 downto 0);
    signal call_457 : std_logic_vector(7 downto 0);
    signal callx_xi363_1500 : std_logic_vector(7 downto 0);
    signal callx_xi_1027 : std_logic_vector(7 downto 0);
    signal cmp161383_1151 : std_logic_vector(0 downto 0);
    signal cmp387_684 : std_logic_vector(0 downto 0);
    signal cmpx_xi368_1524 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1051 : std_logic_vector(0 downto 0);
    signal conv101_815 : std_logic_vector(63 downto 0);
    signal conv107_833 : std_logic_vector(63 downto 0);
    signal conv113_851 : std_logic_vector(63 downto 0);
    signal conv119_869 : std_logic_vector(63 downto 0);
    signal conv125_887 : std_logic_vector(63 downto 0);
    signal conv12_499 : std_logic_vector(15 downto 0);
    signal conv131_905 : std_logic_vector(63 downto 0);
    signal conv145_1103 : std_logic_vector(63 downto 0);
    signal conv147_1107 : std_logic_vector(63 downto 0);
    signal conv150_1111 : std_logic_vector(63 downto 0);
    signal conv153_1115 : std_logic_vector(63 downto 0);
    signal conv155_1145 : std_logic_vector(63 downto 0);
    signal conv165_1253 : std_logic_vector(63 downto 0);
    signal conv170_1266 : std_logic_vector(63 downto 0);
    signal conv176_1284 : std_logic_vector(63 downto 0);
    signal conv182_1302 : std_logic_vector(63 downto 0);
    signal conv188_1320 : std_logic_vector(63 downto 0);
    signal conv194_1338 : std_logic_vector(63 downto 0);
    signal conv19_511 : std_logic_vector(15 downto 0);
    signal conv1_461 : std_logic_vector(31 downto 0);
    signal conv200_1356 : std_logic_vector(63 downto 0);
    signal conv206_1374 : std_logic_vector(63 downto 0);
    signal conv22_524 : std_logic_vector(15 downto 0);
    signal conv230_1715 : std_logic_vector(63 downto 0);
    signal conv255_1671 : std_logic_vector(63 downto 0);
    signal conv261_1675 : std_logic_vector(63 downto 0);
    signal conv263_1664 : std_logic_vector(7 downto 0);
    signal conv289_1723 : std_logic_vector(63 downto 0);
    signal conv297_1732 : std_logic_vector(7 downto 0);
    signal conv29_536 : std_logic_vector(15 downto 0);
    signal conv2x_xi358_1462 : std_logic_vector(31 downto 0);
    signal conv2x_xi_989 : std_logic_vector(31 downto 0);
    signal conv303_1742 : std_logic_vector(7 downto 0);
    signal conv309_1752 : std_logic_vector(7 downto 0);
    signal conv315_1762 : std_logic_vector(7 downto 0);
    signal conv321_1772 : std_logic_vector(7 downto 0);
    signal conv327_1782 : std_logic_vector(7 downto 0);
    signal conv32_549 : std_logic_vector(15 downto 0);
    signal conv333_1792 : std_logic_vector(7 downto 0);
    signal conv339_1802 : std_logic_vector(7 downto 0);
    signal conv39_561 : std_logic_vector(15 downto 0);
    signal conv3_474 : std_logic_vector(31 downto 0);
    signal conv42_574 : std_logic_vector(15 downto 0);
    signal conv49_586 : std_logic_vector(15 downto 0);
    signal conv52_599 : std_logic_vector(15 downto 0);
    signal conv59_611 : std_logic_vector(15 downto 0);
    signal conv5x_xi364_1504 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1031 : std_logic_vector(63 downto 0);
    signal conv62_624 : std_logic_vector(15 downto 0);
    signal conv69_636 : std_logic_vector(15 downto 0);
    signal conv72_649 : std_logic_vector(15 downto 0);
    signal conv79_658 : std_logic_vector(31 downto 0);
    signal conv81_662 : std_logic_vector(31 downto 0);
    signal conv83_678 : std_logic_vector(63 downto 0);
    signal conv90_784 : std_logic_vector(63 downto 0);
    signal conv95_797 : std_logic_vector(63 downto 0);
    signal conv9_486 : std_logic_vector(15 downto 0);
    signal convx_xi367_1519 : std_logic_vector(31 downto 0);
    signal convx_xi_1046 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi362_1478 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_1005 : std_logic_vector(63 downto 0);
    signal exitcond33_925 : std_logic_vector(0 downto 0);
    signal exitcond5_1703 : std_logic_vector(0 downto 0);
    signal exitcond_1394 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1024 : std_logic_vector(15 downto 0);
    signal iNsTr_55_1458 : std_logic_vector(63 downto 0);
    signal iNsTr_65_1497 : std_logic_vector(15 downto 0);
    signal iNsTr_87_1542 : std_logic_vector(63 downto 0);
    signal indvar417_1232 : std_logic_vector(63 downto 0);
    signal indvar431_763 : std_logic_vector(63 downto 0);
    signal indvar_1643 : std_logic_vector(31 downto 0);
    signal indvarx_xnext418_1389 : std_logic_vector(63 downto 0);
    signal indvarx_xnext432_920 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1698 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_957 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1426 : std_logic_vector(63 downto 0);
    signal mul148_1120 : std_logic_vector(63 downto 0);
    signal mul151_1125 : std_logic_vector(63 downto 0);
    signal mul154_1130 : std_logic_vector(63 downto 0);
    signal mul236_1581 : std_logic_vector(15 downto 0);
    signal mul249_1594 : std_logic_vector(15 downto 0);
    signal mul254_1655 : std_logic_vector(31 downto 0);
    signal mul260_1660 : std_logic_vector(31 downto 0);
    signal mul82_672 : std_logic_vector(31 downto 0);
    signal mul_667 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi361_1471 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_998 : std_logic_vector(15 downto 0);
    signal phitmp391_1423 : std_logic_vector(63 downto 0);
    signal phitmp_954 : std_logic_vector(63 downto 0);
    signal ptr_deref_1095_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1095_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1095_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1095_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1095_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1095_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1381_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1381_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1381_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1381_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1381_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1381_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1568_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1568_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1568_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1568_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1568_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1568_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_912_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_912_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_912_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_912_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_912_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_912_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1136 : std_logic_vector(63 downto 0);
    signal sh_promx_xi375_1554 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1081 : std_logic_vector(63 downto 0);
    signal shl104_826 : std_logic_vector(63 downto 0);
    signal shl10_492 : std_logic_vector(15 downto 0);
    signal shl110_844 : std_logic_vector(63 downto 0);
    signal shl116_862 : std_logic_vector(63 downto 0);
    signal shl122_880 : std_logic_vector(63 downto 0);
    signal shl128_898 : std_logic_vector(63 downto 0);
    signal shl14x_xi376_1559 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1086 : std_logic_vector(63 downto 0);
    signal shl167_1259 : std_logic_vector(63 downto 0);
    signal shl173_1277 : std_logic_vector(63 downto 0);
    signal shl179_1295 : std_logic_vector(63 downto 0);
    signal shl185_1313 : std_logic_vector(63 downto 0);
    signal shl191_1331 : std_logic_vector(63 downto 0);
    signal shl197_1349 : std_logic_vector(63 downto 0);
    signal shl203_1367 : std_logic_vector(63 downto 0);
    signal shl20_517 : std_logic_vector(15 downto 0);
    signal shl30_542 : std_logic_vector(15 downto 0);
    signal shl40_567 : std_logic_vector(15 downto 0);
    signal shl50_592 : std_logic_vector(15 downto 0);
    signal shl60_617 : std_logic_vector(15 downto 0);
    signal shl70_642 : std_logic_vector(15 downto 0);
    signal shl8x_xi366_1515 : std_logic_vector(63 downto 0);
    signal shl8x_xi366x_xlcssa_1532 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1042 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1059 : std_logic_vector(63 downto 0);
    signal shl92_790 : std_logic_vector(63 downto 0);
    signal shl98_808 : std_logic_vector(63 downto 0);
    signal shl_467 : std_logic_vector(31 downto 0);
    signal shlx_xi359_1468 : std_logic_vector(31 downto 0);
    signal shlx_xi_995 : std_logic_vector(31 downto 0);
    signal shr300_1738 : std_logic_vector(63 downto 0);
    signal shr306_1748 : std_logic_vector(63 downto 0);
    signal shr312_1758 : std_logic_vector(63 downto 0);
    signal shr318_1768 : std_logic_vector(63 downto 0);
    signal shr324_1778 : std_logic_vector(63 downto 0);
    signal shr330_1788 : std_logic_vector(63 downto 0);
    signal shr336_1798 : std_logic_vector(63 downto 0);
    signal sub273_1606 : std_logic_vector(15 downto 0);
    signal sub293_1728 : std_logic_vector(63 downto 0);
    signal sub_1600 : std_logic_vector(15 downto 0);
    signal tmp13_1174 : std_logic_vector(63 downto 0);
    signal tmp14_1178 : std_logic_vector(63 downto 0);
    signal tmp15_1183 : std_logic_vector(63 downto 0);
    signal tmp16_1187 : std_logic_vector(63 downto 0);
    signal tmp17_1192 : std_logic_vector(63 downto 0);
    signal tmp18_1196 : std_logic_vector(63 downto 0);
    signal tmp19_1201 : std_logic_vector(63 downto 0);
    signal tmp20_1205 : std_logic_vector(31 downto 0);
    signal tmp21_1210 : std_logic_vector(63 downto 0);
    signal tmp22_1216 : std_logic_vector(63 downto 0);
    signal tmp23_1222 : std_logic_vector(0 downto 0);
    signal tmp25_722 : std_logic_vector(31 downto 0);
    signal tmp26_727 : std_logic_vector(31 downto 0);
    signal tmp27_731 : std_logic_vector(31 downto 0);
    signal tmp28_736 : std_logic_vector(31 downto 0);
    signal tmp29_741 : std_logic_vector(63 downto 0);
    signal tmp30_747 : std_logic_vector(63 downto 0);
    signal tmp31_753 : std_logic_vector(0 downto 0);
    signal tmp392_1491 : std_logic_vector(15 downto 0);
    signal tmp393_1612 : std_logic_vector(15 downto 0);
    signal tmp3_1616 : std_logic_vector(31 downto 0);
    signal tmp412_1164 : std_logic_vector(63 downto 0);
    signal tmp413_1170 : std_logic_vector(0 downto 0);
    signal tmp414_1414 : std_logic_vector(63 downto 0);
    signal tmp421_696 : std_logic_vector(31 downto 0);
    signal tmp423_701 : std_logic_vector(31 downto 0);
    signal tmp424_706 : std_logic_vector(63 downto 0);
    signal tmp425_712 : std_logic_vector(63 downto 0);
    signal tmp426_718 : std_logic_vector(0 downto 0);
    signal tmp428_945 : std_logic_vector(63 downto 0);
    signal tmp4_1622 : std_logic_vector(31 downto 0);
    signal tmp6_1626 : std_logic_vector(31 downto 0);
    signal tmp7_1631 : std_logic_vector(15 downto 0);
    signal tmp8_1635 : std_logic_vector(31 downto 0);
    signal tmp9_1640 : std_logic_vector(31 downto 0);
    signal tmp_1018 : std_logic_vector(15 downto 0);
    signal tobool218_1445 : std_logic_vector(0 downto 0);
    signal tobool_976 : std_logic_vector(0 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1004_wire : std_logic_vector(15 downto 0);
    signal type_cast_1009_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1011_wire : std_logic_vector(63 downto 0);
    signal type_cast_1016_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1022_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1040_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1062_wire : std_logic_vector(63 downto 0);
    signal type_cast_1067_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1073_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1079_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1139_wire : std_logic_vector(63 downto 0);
    signal type_cast_1142_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1162_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1208_wire : std_logic_vector(63 downto 0);
    signal type_cast_1214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1220_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1238_wire : std_logic_vector(63 downto 0);
    signal type_cast_1257_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1275_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1311_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1329_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1347_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1365_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1387_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1417_wire : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1429_wire : std_logic_vector(63 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1466_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1477_wire : std_logic_vector(15 downto 0);
    signal type_cast_1482_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1484_wire : std_logic_vector(63 downto 0);
    signal type_cast_1489_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1495_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1535_wire : std_logic_vector(63 downto 0);
    signal type_cast_1540_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1546_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1552_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1598_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1610_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1646_wire : std_logic_vector(31 downto 0);
    signal type_cast_1649_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1679_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1713_wire : std_logic_vector(63 downto 0);
    signal type_cast_1721_wire : std_logic_vector(63 downto 0);
    signal type_cast_1736_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1746_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1766_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1776_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1786_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_465_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_490_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_515_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_540_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_615_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_640_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_676_wire : std_logic_vector(63 downto 0);
    signal type_cast_682_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_704_wire : std_logic_vector(63 downto 0);
    signal type_cast_710_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_739_wire : std_logic_vector(63 downto 0);
    signal type_cast_745_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_751_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_758_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_766_wire : std_logic_vector(63 downto 0);
    signal type_cast_769_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_806_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_842_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_860_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_896_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_918_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_937_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire : std_logic_vector(63 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_960_wire : std_logic_vector(63 downto 0);
    signal type_cast_963_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_968_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_974_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_987_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_993_wire_constant : std_logic_vector(31 downto 0);
    signal umax24_1229 : std_logic_vector(63 downto 0);
    signal umax32_760 : std_logic_vector(63 downto 0);
    signal umax427_939 : std_logic_vector(63 downto 0);
    signal umax_1408 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1091_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1091_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1091_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1091_resized_base_address <= "00000000000000";
    array_obj_ref_1244_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1244_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1244_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1244_resized_base_address <= "00000000000000";
    array_obj_ref_1564_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1564_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1564_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1564_resized_base_address <= "00000000000000";
    array_obj_ref_775_constant_part_of_offset <= "00000000000000";
    array_obj_ref_775_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_775_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_775_resized_base_address <= "00000000000000";
    ptr_deref_1095_word_offset_0 <= "00000000000000";
    ptr_deref_1381_word_offset_0 <= "00000000000000";
    ptr_deref_1568_word_offset_0 <= "00000000000000";
    ptr_deref_912_word_offset_0 <= "00000000000000";
    type_cast_1002_wire_constant <= "0000000000000000";
    type_cast_1009_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1016_wire_constant <= "0000000000000001";
    type_cast_1022_wire_constant <= "0000000000000001";
    type_cast_1040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1067_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1073_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1079_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1134_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1142_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1149_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1162_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1168_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1220_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1227_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1257_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1275_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1293_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1329_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1347_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1365_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1387_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1406_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1432_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1456_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1466_wire_constant <= "00000000000000000000000000000110";
    type_cast_1475_wire_constant <= "0000000000000000";
    type_cast_1482_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1489_wire_constant <= "0000000000000001";
    type_cast_1495_wire_constant <= "0000000000000001";
    type_cast_1513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1540_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1546_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1552_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1584_wire_constant <= "11001000";
    type_cast_1588_wire_constant <= "11001000";
    type_cast_1598_wire_constant <= "1111111111111111";
    type_cast_1604_wire_constant <= "1111111111111111";
    type_cast_1610_wire_constant <= "1111111111111111";
    type_cast_1620_wire_constant <= "00000000000000000000000000000001";
    type_cast_1649_wire_constant <= "00000000000000000000000000000000";
    type_cast_1679_wire_constant <= "00000001";
    type_cast_1696_wire_constant <= "00000000000000000000000000000001";
    type_cast_1736_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1746_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1766_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1776_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1786_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_465_wire_constant <= "00000000000000000000000000001000";
    type_cast_490_wire_constant <= "0000000000001000";
    type_cast_515_wire_constant <= "0000000000001000";
    type_cast_540_wire_constant <= "0000000000001000";
    type_cast_565_wire_constant <= "0000000000001000";
    type_cast_590_wire_constant <= "0000000000001000";
    type_cast_615_wire_constant <= "0000000000001000";
    type_cast_640_wire_constant <= "0000000000001000";
    type_cast_682_wire_constant <= "00000000000000000000000000000011";
    type_cast_710_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_745_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_751_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_758_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_769_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_806_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_824_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_860_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_878_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_896_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_918_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_937_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_951_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_963_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_968_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_974_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_987_wire_constant <= "00000000000000000000000000000001";
    type_cast_993_wire_constant <= "00000000000000000000000000000110";
    phi_stmt_1005: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1009_wire_constant & type_cast_1011_wire;
      req <= phi_stmt_1005_req_0 & phi_stmt_1005_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1005",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1005_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_1005,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1005
    phi_stmt_1059: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1062_wire;
      req(0) <= phi_stmt_1059_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1059",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1059_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1059
    phi_stmt_1232: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1236_wire_constant & type_cast_1238_wire;
      req <= phi_stmt_1232_req_0 & phi_stmt_1232_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1232",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1232_ack_0,
          idata => idata,
          odata => indvar417_1232,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1232
    phi_stmt_1426: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1429_wire & type_cast_1432_wire_constant;
      req <= phi_stmt_1426_req_0 & phi_stmt_1426_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1426",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1426_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1426,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1426
    phi_stmt_1471: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1475_wire_constant & type_cast_1477_wire;
      req <= phi_stmt_1471_req_0 & phi_stmt_1471_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1471",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1471_ack_0,
          idata => idata,
          odata => nx_x022x_xi361_1471,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1471
    phi_stmt_1478: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1482_wire_constant & type_cast_1484_wire;
      req <= phi_stmt_1478_req_0 & phi_stmt_1478_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1478",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1478_ack_0,
          idata => idata,
          odata => elementx_x021x_xi362_1478,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1478
    phi_stmt_1532: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1535_wire;
      req(0) <= phi_stmt_1532_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1532",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1532_ack_0,
          idata => idata,
          odata => shl8x_xi366x_xlcssa_1532,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1532
    phi_stmt_1643: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1646_wire & type_cast_1649_wire_constant;
      req <= phi_stmt_1643_req_0 & phi_stmt_1643_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1643",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1643_ack_0,
          idata => idata,
          odata => indvar_1643,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1643
    phi_stmt_763: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_766_wire & type_cast_769_wire_constant;
      req <= phi_stmt_763_req_0 & phi_stmt_763_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_763",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_763_ack_0,
          idata => idata,
          odata => indvar431_763,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_763
    phi_stmt_957: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_960_wire & type_cast_963_wire_constant;
      req <= phi_stmt_957_req_0 & phi_stmt_957_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_957",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_957_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_957,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_957
    phi_stmt_998: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1002_wire_constant & type_cast_1004_wire;
      req <= phi_stmt_998_req_0 & phi_stmt_998_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_998",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_998_ack_0,
          idata => idata,
          odata => nx_x022x_xi_998,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_998
    -- flow-through select operator MUX_1228_inst
    umax24_1229 <= tmp22_1216 when (tmp23_1222(0) /=  '0') else type_cast_1227_wire_constant;
    -- flow-through select operator MUX_1407_inst
    umax_1408 <= tmp412_1164 when (tmp413_1170(0) /=  '0') else type_cast_1406_wire_constant;
    -- flow-through select operator MUX_759_inst
    umax32_760 <= tmp30_747 when (tmp31_753(0) /=  '0') else type_cast_758_wire_constant;
    -- flow-through select operator MUX_938_inst
    umax427_939 <= tmp425_712 when (tmp426_718(0) /=  '0') else type_cast_937_wire_constant;
    addr_of_1092_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1092_final_reg_req_0;
      addr_of_1092_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1092_final_reg_req_1;
      addr_of_1092_final_reg_ack_1<= rack(0);
      addr_of_1092_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1092_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1091_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1245_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1245_final_reg_req_0;
      addr_of_1245_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1245_final_reg_req_1;
      addr_of_1245_final_reg_ack_1<= rack(0);
      addr_of_1245_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1245_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1244_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1565_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1565_final_reg_req_0;
      addr_of_1565_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1565_final_reg_req_1;
      addr_of_1565_final_reg_ack_1<= rack(0);
      addr_of_1565_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1565_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1564_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1566,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_776_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_776_final_reg_req_0;
      addr_of_776_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_776_final_reg_req_1;
      addr_of_776_final_reg_ack_1<= rack(0);
      addr_of_776_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_776_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_775_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1004_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1004_inst_req_0;
      type_cast_1004_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1004_inst_req_1;
      type_cast_1004_inst_ack_1<= rack(0);
      type_cast_1004_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1004_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1024,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1004_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1011_inst_req_0;
      type_cast_1011_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1011_inst_req_1;
      type_cast_1011_inst_ack_1<= rack(0);
      type_cast_1011_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1042,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1011_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1030_inst_req_0;
      type_cast_1030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1030_inst_req_1;
      type_cast_1030_inst_ack_1<= rack(0);
      type_cast_1030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1045_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1045_inst_req_0;
      type_cast_1045_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1045_inst_req_1;
      type_cast_1045_inst_ack_1<= rack(0);
      type_cast_1045_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1045_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1046,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1062_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1062_inst_req_0;
      type_cast_1062_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1062_inst_req_1;
      type_cast_1062_inst_ack_1<= rack(0);
      type_cast_1062_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1062_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1042,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1062_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1102_inst_req_0;
      type_cast_1102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1102_inst_req_1;
      type_cast_1102_inst_ack_1<= rack(0);
      type_cast_1102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1114_inst_req_0;
      type_cast_1114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1114_inst_req_1;
      type_cast_1114_inst_ack_1<= rack(0);
      type_cast_1114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1139_inst
    process(sext_1136) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1136(63 downto 0);
      type_cast_1139_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1144_inst
    process(ASHR_i64_i64_1143_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1143_wire(63 downto 0);
      conv155_1145 <= tmp_var; -- 
    end process;
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1177_inst_req_0;
      type_cast_1177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1177_inst_req_1;
      type_cast_1177_inst_ack_1<= rack(0);
      type_cast_1177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp14_1178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1186_inst_req_0;
      type_cast_1186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1186_inst_req_1;
      type_cast_1186_inst_ack_1<= rack(0);
      type_cast_1186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_1187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1195_inst_req_0;
      type_cast_1195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1195_inst_req_1;
      type_cast_1195_inst_ack_1<= rack(0);
      type_cast_1195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_654,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp18_1196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1204_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1204_inst_req_0;
      type_cast_1204_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1204_inst_req_1;
      type_cast_1204_inst_ack_1<= rack(0);
      type_cast_1204_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1204_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp19_1201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1209_inst_req_0;
      type_cast_1209_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1209_inst_req_1;
      type_cast_1209_inst_ack_1<= rack(0);
      type_cast_1209_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1208_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp21_1210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext418_1389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1238_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1252_inst_req_0;
      type_cast_1252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1252_inst_req_1;
      type_cast_1252_inst_ack_1<= rack(0);
      type_cast_1252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1249,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1265_inst_req_0;
      type_cast_1265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1265_inst_req_1;
      type_cast_1265_inst_ack_1<= rack(0);
      type_cast_1265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1283_inst_req_0;
      type_cast_1283_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1283_inst_req_1;
      type_cast_1283_inst_ack_1<= rack(0);
      type_cast_1283_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1283_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1284,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1301_inst_req_0;
      type_cast_1301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1301_inst_req_1;
      type_cast_1301_inst_ack_1<= rack(0);
      type_cast_1301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1319_inst_req_0;
      type_cast_1319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1319_inst_req_1;
      type_cast_1319_inst_ack_1<= rack(0);
      type_cast_1319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1337_inst_req_0;
      type_cast_1337_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1337_inst_req_1;
      type_cast_1337_inst_ack_1<= rack(0);
      type_cast_1337_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1337_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1334,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1338,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1355_inst_req_0;
      type_cast_1355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1355_inst_req_1;
      type_cast_1355_inst_ack_1<= rack(0);
      type_cast_1355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1373_inst_req_0;
      type_cast_1373_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1373_inst_req_1;
      type_cast_1373_inst_ack_1<= rack(0);
      type_cast_1373_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1373_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1374,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1417_inst
    process(tmp414_1414) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp414_1414(63 downto 0);
      type_cast_1417_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1422_inst
    process(ASHR_i64_i64_1421_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1421_wire(63 downto 0);
      phitmp391_1423 <= tmp_var; -- 
    end process;
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp391_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1429_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1461_inst_req_0;
      type_cast_1461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1461_inst_req_1;
      type_cast_1461_inst_ack_1<= rack(0);
      type_cast_1461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_55_1458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi358_1462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1477_inst_req_0;
      type_cast_1477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1477_inst_req_1;
      type_cast_1477_inst_ack_1<= rack(0);
      type_cast_1477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_65_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1477_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1484_inst_req_0;
      type_cast_1484_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1484_inst_req_1;
      type_cast_1484_inst_ack_1<= rack(0);
      type_cast_1484_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1484_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi366_1515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1484_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1503_inst_req_0;
      type_cast_1503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1503_inst_req_1;
      type_cast_1503_inst_ack_1<= rack(0);
      type_cast_1503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi363_1500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi364_1504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1518_inst_req_0;
      type_cast_1518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1518_inst_req_1;
      type_cast_1518_inst_ack_1<= rack(0);
      type_cast_1518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp392_1491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi367_1519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1535_inst_req_0;
      type_cast_1535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1535_inst_req_1;
      type_cast_1535_inst_ack_1<= rack(0);
      type_cast_1535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi366_1515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1535_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1615_inst_req_0;
      type_cast_1615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1615_inst_req_1;
      type_cast_1615_inst_ack_1<= rack(0);
      type_cast_1615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp393_1612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1634_inst_req_0;
      type_cast_1634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1634_inst_req_1;
      type_cast_1634_inst_ack_1<= rack(0);
      type_cast_1634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1646_inst_req_0;
      type_cast_1646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1646_inst_req_1;
      type_cast_1646_inst_ack_1<= rack(0);
      type_cast_1646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1646_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1663_inst_req_0;
      type_cast_1663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1663_inst_req_1;
      type_cast_1663_inst_ack_1<= rack(0);
      type_cast_1663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvar_1643,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1670_inst_req_0;
      type_cast_1670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1670_inst_req_1;
      type_cast_1670_inst_ack_1<= rack(0);
      type_cast_1670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul254_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1674_inst_req_0;
      type_cast_1674_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1674_inst_req_1;
      type_cast_1674_inst_ack_1<= rack(0);
      type_cast_1674_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1674_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul260_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv261_1675,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1714_inst_req_0;
      type_cast_1714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1714_inst_req_1;
      type_cast_1714_inst_ack_1<= rack(0);
      type_cast_1714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1713_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1722_inst_req_0;
      type_cast_1722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1722_inst_req_1;
      type_cast_1722_inst_ack_1<= rack(0);
      type_cast_1722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1721_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv289_1723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1731_inst_req_0;
      type_cast_1731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1731_inst_req_1;
      type_cast_1731_inst_ack_1<= rack(0);
      type_cast_1731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub293_1728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv297_1732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1741_inst_req_0;
      type_cast_1741_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1741_inst_req_1;
      type_cast_1741_inst_ack_1<= rack(0);
      type_cast_1741_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1741_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr300_1738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv303_1742,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1751_inst_req_0;
      type_cast_1751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1751_inst_req_1;
      type_cast_1751_inst_ack_1<= rack(0);
      type_cast_1751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr306_1748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv309_1752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1761_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1761_inst_req_0;
      type_cast_1761_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1761_inst_req_1;
      type_cast_1761_inst_ack_1<= rack(0);
      type_cast_1761_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1761_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr312_1758,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv315_1762,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1771_inst_req_0;
      type_cast_1771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1771_inst_req_1;
      type_cast_1771_inst_ack_1<= rack(0);
      type_cast_1771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1771_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr318_1768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv321_1772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1781_inst_req_0;
      type_cast_1781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1781_inst_req_1;
      type_cast_1781_inst_ack_1<= rack(0);
      type_cast_1781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr324_1778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv327_1782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1791_inst_req_0;
      type_cast_1791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1791_inst_req_1;
      type_cast_1791_inst_ack_1<= rack(0);
      type_cast_1791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr330_1788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv333_1792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1801_inst_req_0;
      type_cast_1801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1801_inst_req_1;
      type_cast_1801_inst_ack_1<= rack(0);
      type_cast_1801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr336_1798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_460_inst_req_0;
      type_cast_460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_460_inst_req_1;
      type_cast_460_inst_ack_1<= rack(0);
      type_cast_460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_498_inst_req_0;
      type_cast_498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_498_inst_req_1;
      type_cast_498_inst_ack_1<= rack(0);
      type_cast_498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_510_inst_req_0;
      type_cast_510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_510_inst_req_1;
      type_cast_510_inst_ack_1<= rack(0);
      type_cast_510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_511,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_523_inst_req_0;
      type_cast_523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_523_inst_req_1;
      type_cast_523_inst_ack_1<= rack(0);
      type_cast_523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_535_inst_req_0;
      type_cast_535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_535_inst_req_1;
      type_cast_535_inst_ack_1<= rack(0);
      type_cast_535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_532,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_548_inst_req_0;
      type_cast_548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_548_inst_req_1;
      type_cast_548_inst_ack_1<= rack(0);
      type_cast_548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_560_inst_req_0;
      type_cast_560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_560_inst_req_1;
      type_cast_560_inst_ack_1<= rack(0);
      type_cast_560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_573_inst_req_0;
      type_cast_573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_573_inst_req_1;
      type_cast_573_inst_ack_1<= rack(0);
      type_cast_573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_585_inst_req_0;
      type_cast_585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_585_inst_req_1;
      type_cast_585_inst_ack_1<= rack(0);
      type_cast_585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_582,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_635_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_635_inst_req_0;
      type_cast_635_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_635_inst_req_1;
      type_cast_635_inst_ack_1<= rack(0);
      type_cast_635_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_635_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_632,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_648_inst_req_0;
      type_cast_648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_648_inst_req_1;
      type_cast_648_inst_ack_1<= rack(0);
      type_cast_648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_657_inst_req_0;
      type_cast_657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_657_inst_req_1;
      type_cast_657_inst_ack_1<= rack(0);
      type_cast_657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_661_inst_req_0;
      type_cast_661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_661_inst_req_1;
      type_cast_661_inst_ack_1<= rack(0);
      type_cast_661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_677_inst_req_0;
      type_cast_677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_677_inst_req_1;
      type_cast_677_inst_ack_1<= rack(0);
      type_cast_677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_676_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_705_inst_req_0;
      type_cast_705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_705_inst_req_1;
      type_cast_705_inst_ack_1<= rack(0);
      type_cast_705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_704_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp424_706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_721_inst_req_0;
      type_cast_721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_721_inst_req_1;
      type_cast_721_inst_ack_1<= rack(0);
      type_cast_721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp25_722,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_730_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_730_inst_req_0;
      type_cast_730_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_730_inst_req_1;
      type_cast_730_inst_ack_1<= rack(0);
      type_cast_730_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_730_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp27_731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_740_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_740_inst_req_0;
      type_cast_740_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_740_inst_req_1;
      type_cast_740_inst_ack_1<= rack(0);
      type_cast_740_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_740_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_739_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp29_741,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_766_inst_req_0;
      type_cast_766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_766_inst_req_1;
      type_cast_766_inst_ack_1<= rack(0);
      type_cast_766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext432_920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_766_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_783_inst_req_0;
      type_cast_783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_783_inst_req_1;
      type_cast_783_inst_ack_1<= rack(0);
      type_cast_783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_796_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_796_inst_req_0;
      type_cast_796_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_796_inst_req_1;
      type_cast_796_inst_ack_1<= rack(0);
      type_cast_796_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_796_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_829,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_850_inst_req_0;
      type_cast_850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_850_inst_req_1;
      type_cast_850_inst_ack_1<= rack(0);
      type_cast_850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_868_inst_req_0;
      type_cast_868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_868_inst_req_1;
      type_cast_868_inst_ack_1<= rack(0);
      type_cast_868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_865,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_869,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_886_inst_req_0;
      type_cast_886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_886_inst_req_1;
      type_cast_886_inst_ack_1<= rack(0);
      type_cast_886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_904_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_904_inst_req_0;
      type_cast_904_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_904_inst_req_1;
      type_cast_904_inst_ack_1<= rack(0);
      type_cast_904_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_904_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_901,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_905,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_948_inst
    process(tmp428_945) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp428_945(63 downto 0);
      type_cast_948_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_953_inst
    process(ASHR_i64_i64_952_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_952_wire(63 downto 0);
      phitmp_954 <= tmp_var; -- 
    end process;
    type_cast_960_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_960_inst_req_0;
      type_cast_960_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_960_inst_req_1;
      type_cast_960_inst_ack_1<= rack(0);
      type_cast_960_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_960_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_954,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_960_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1091_index_1_rename
    process(R_ix_x0x_xlcssa_1090_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1090_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1090_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1091_index_1_resize
    process(ix_x0x_xlcssa_957) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_957;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1090_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1091_root_address_inst
    process(array_obj_ref_1091_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1091_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1091_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_index_1_rename
    process(R_indvar417_1243_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar417_1243_resized;
      ov(13 downto 0) := iv;
      R_indvar417_1243_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_index_1_resize
    process(indvar417_1232) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar417_1232;
      ov := iv(13 downto 0);
      R_indvar417_1243_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1244_root_address_inst
    process(array_obj_ref_1244_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1244_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1244_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1564_index_1_rename
    process(R_ix_x1x_xlcssa_1563_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1563_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1563_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1564_index_1_resize
    process(ix_x1x_xlcssa_1426) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1426;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1563_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1564_root_address_inst
    process(array_obj_ref_1564_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1564_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1564_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_775_index_1_rename
    process(R_indvar431_774_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar431_774_resized;
      ov(13 downto 0) := iv;
      R_indvar431_774_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_775_index_1_resize
    process(indvar431_763) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar431_763;
      ov := iv(13 downto 0);
      R_indvar431_774_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_775_root_address_inst
    process(array_obj_ref_775_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_775_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_775_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1095_addr_0
    process(ptr_deref_1095_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1095_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1095_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1095_base_resize
    process(arrayidx143_1093) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1093;
      ov := iv(13 downto 0);
      ptr_deref_1095_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1095_gather_scatter
    process(shl14x_xi_1086) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1086;
      ov(63 downto 0) := iv;
      ptr_deref_1095_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1095_root_address_inst
    process(ptr_deref_1095_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1095_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1095_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1381_addr_0
    process(ptr_deref_1381_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1381_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1381_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1381_base_resize
    process(arrayidx211_1246) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1246;
      ov := iv(13 downto 0);
      ptr_deref_1381_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1381_gather_scatter
    process(add207_1379) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1379;
      ov(63 downto 0) := iv;
      ptr_deref_1381_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1381_root_address_inst
    process(ptr_deref_1381_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1381_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1381_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1568_addr_0
    process(ptr_deref_1568_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1568_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1568_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1568_base_resize
    process(arrayidx226_1566) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1566;
      ov := iv(13 downto 0);
      ptr_deref_1568_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1568_gather_scatter
    process(shl14x_xi376_1559) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi376_1559;
      ov(63 downto 0) := iv;
      ptr_deref_1568_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1568_root_address_inst
    process(ptr_deref_1568_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1568_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1568_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_912_addr_0
    process(ptr_deref_912_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_912_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_912_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_912_base_resize
    process(arrayidx_777) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_777;
      ov := iv(13 downto 0);
      ptr_deref_912_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_912_gather_scatter
    process(add132_910) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_910;
      ov(63 downto 0) := iv;
      ptr_deref_912_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_912_root_address_inst
    process(ptr_deref_912_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_912_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_912_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1052_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1051;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1052_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1052_branch_req_0,
          ack0 => if_stmt_1052_branch_ack_0,
          ack1 => if_stmt_1052_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1152_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161383_1151;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1152_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1152_branch_req_0,
          ack0 => if_stmt_1152_branch_ack_0,
          ack1 => if_stmt_1152_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1395_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1394;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1395_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1395_branch_req_0,
          ack0 => if_stmt_1395_branch_ack_0,
          ack1 => if_stmt_1395_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1446_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1445;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1446_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1446_branch_req_0,
          ack0 => if_stmt_1446_branch_ack_0,
          ack1 => if_stmt_1446_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1525_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi368_1524;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1525_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1525_branch_req_0,
          ack0 => if_stmt_1525_branch_ack_0,
          ack1 => if_stmt_1525_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1704_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1703;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1704_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1704_branch_req_0,
          ack0 => if_stmt_1704_branch_ack_0,
          ack1 => if_stmt_1704_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_685_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp387_684;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_685_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_685_branch_req_0,
          ack0 => if_stmt_685_branch_ack_0,
          ack1 => if_stmt_685_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_926_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond33_925;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_926_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_926_branch_req_0,
          ack0 => if_stmt_926_branch_ack_0,
          ack1 => if_stmt_926_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_977_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_976;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_977_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_977_branch_req_0,
          ack0 => if_stmt_977_branch_ack_0,
          ack1 => if_stmt_977_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1017_inst
    process(nx_x022x_xi_998) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_998, type_cast_1016_wire_constant, tmp_var);
      tmp_1018 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1023_inst
    process(nx_x022x_xi_998) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_998, type_cast_1022_wire_constant, tmp_var);
      iNsTr_35_1024 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1490_inst
    process(nx_x022x_xi361_1471) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi361_1471, type_cast_1489_wire_constant, tmp_var);
      tmp392_1491 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1496_inst
    process(nx_x022x_xi361_1471) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi361_1471, type_cast_1495_wire_constant, tmp_var);
      iNsTr_65_1497 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1599_inst
    process(add43_579) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43_579, type_cast_1598_wire_constant, tmp_var);
      sub_1600 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1605_inst
    process(add63_629) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add63_629, type_cast_1604_wire_constant, tmp_var);
      sub273_1606 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1611_inst
    process(add53_604) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_604, type_cast_1610_wire_constant, tmp_var);
      tmp393_1612 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1621_inst
    process(tmp3_1616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1616, type_cast_1620_wire_constant, tmp_var);
      tmp4_1622 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1659_inst
    process(tmp9_1640, mul254_1655) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1640, mul254_1655, tmp_var);
      mul260_1660 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1697_inst
    process(indvar_1643) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1643, type_cast_1696_wire_constant, tmp_var);
      indvarx_xnext_1698 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1388_inst
    process(indvar417_1232) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar417_1232, type_cast_1387_wire_constant, tmp_var);
      indvarx_xnext418_1389 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_919_inst
    process(indvar431_763) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar431_763, type_cast_918_wire_constant, tmp_var);
      indvarx_xnext432_920 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1467_inst
    process(conv2x_xi358_1462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi358_1462, type_cast_1466_wire_constant, tmp_var);
      shlx_xi359_1468 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_994_inst
    process(conv2x_xi_989) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_989, type_cast_993_wire_constant, tmp_var);
      shlx_xi_995 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1074_inst
    process(Bx_xnot_1069) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1069, type_cast_1073_wire_constant, tmp_var);
      add1216x_xi_1075 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1438_inst
    process(conv155_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1145, type_cast_1437_wire_constant, tmp_var);
      and217_1439 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1547_inst
    process(iNsTr_87_1542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_87_1542, type_cast_1546_wire_constant, tmp_var);
      add1216x_xi374_1548 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_969_inst
    process(conv83_678) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_678, type_cast_968_wire_constant, tmp_var);
      and_970 <= tmp_var; --
    end process;
    -- binary operator AND_u8_u8_1680_inst
    process(conv263_1664) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv263_1664, type_cast_1679_wire_constant, tmp_var);
      and264_1681 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1143_inst
    process(type_cast_1139_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1139_wire, type_cast_1142_wire_constant, tmp_var);
      ASHR_i64_i64_1143_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1421_inst
    process(type_cast_1417_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1417_wire, type_cast_1420_wire_constant, tmp_var);
      ASHR_i64_i64_1421_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_952_inst
    process(type_cast_948_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_948_wire, type_cast_951_wire_constant, tmp_var);
      ASHR_i64_i64_952_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1702_inst
    process(indvarx_xnext_1698, tmp4_1622) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1698, tmp4_1622, tmp_var);
      exitcond5_1703 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1393_inst
    process(indvarx_xnext418_1389, umax24_1229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext418_1389, umax24_1229, tmp_var);
      exitcond_1394 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1444_inst
    process(and217_1439) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1439, type_cast_1443_wire_constant, tmp_var);
      tobool218_1445 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_924_inst
    process(indvarx_xnext432_920, umax32_760) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext432_920, umax32_760, tmp_var);
      exitcond33_925 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_975_inst
    process(and_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_970, type_cast_974_wire_constant, tmp_var);
      tobool_976 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1163_inst
    process(conv155_1145) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1145, type_cast_1162_wire_constant, tmp_var);
      tmp412_1164 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1215_inst
    process(tmp21_1210) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp21_1210, type_cast_1214_wire_constant, tmp_var);
      tmp22_1216 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1737_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1736_wire_constant, tmp_var);
      shr300_1738 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1747_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1746_wire_constant, tmp_var);
      shr306_1748 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1757_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1756_wire_constant, tmp_var);
      shr312_1758 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1767_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1766_wire_constant, tmp_var);
      shr318_1768 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1777_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1776_wire_constant, tmp_var);
      shr324_1778 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1787_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1786_wire_constant, tmp_var);
      shr330_1788 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1797_inst
    process(sub293_1728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub293_1728, type_cast_1796_wire_constant, tmp_var);
      shr336_1798 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_711_inst
    process(tmp424_706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp424_706, type_cast_710_wire_constant, tmp_var);
      tmp425_712 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_746_inst
    process(tmp29_741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp29_741, type_cast_745_wire_constant, tmp_var);
      tmp30_747 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1580_inst
    process(add73_654, add23_529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_654, add23_529, tmp_var);
      mul236_1581 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1593_inst
    process(add43_579, add33_554) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_579, add33_554, tmp_var);
      mul249_1594 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1630_inst
    process(add73_654, add23_529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_654, add23_529, tmp_var);
      tmp7_1631 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1639_inst
    process(tmp6_1626, tmp8_1635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1626, tmp8_1635, tmp_var);
      tmp9_1640 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1654_inst
    process(tmp9_1640, indvar_1643) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1640, indvar_1643, tmp_var);
      mul254_1655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_666_inst
    process(conv79_658, add_479) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_658, add_479, tmp_var);
      mul_667 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_671_inst
    process(mul_667, conv81_662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_667, conv81_662, tmp_var);
      mul82_672 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_695_inst
    process(add_479, conv79_658) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_479, conv79_658, tmp_var);
      tmp421_696 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_700_inst
    process(tmp421_696, conv81_662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp421_696, conv81_662, tmp_var);
      tmp423_701 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_726_inst
    process(add_479, tmp25_722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_479, tmp25_722, tmp_var);
      tmp26_727 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_735_inst
    process(tmp26_727, tmp27_731) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_727, tmp27_731, tmp_var);
      tmp28_736 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1119_inst
    process(conv153_1115, conv145_1103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1115, conv145_1103, tmp_var);
      mul148_1120 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1124_inst
    process(mul148_1120, conv150_1111) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1120, conv150_1111, tmp_var);
      mul151_1125 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1129_inst
    process(mul151_1125, conv147_1107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1125, conv147_1107, tmp_var);
      mul154_1130 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1182_inst
    process(tmp13_1174, tmp14_1178) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_1174, tmp14_1178, tmp_var);
      tmp15_1183 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1191_inst
    process(tmp15_1183, tmp16_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp15_1183, tmp16_1187, tmp_var);
      tmp17_1192 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1200_inst
    process(tmp17_1192, tmp18_1196) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp17_1192, tmp18_1196, tmp_var);
      tmp19_1201 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_503_inst
    process(shl10_492, conv12_499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_492, conv12_499, tmp_var);
      add13_504 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_528_inst
    process(shl20_517, conv22_524) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_517, conv22_524, tmp_var);
      add23_529 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_553_inst
    process(shl30_542, conv32_549) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_542, conv32_549, tmp_var);
      add33_554 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_578_inst
    process(shl40_567, conv42_574) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_567, conv42_574, tmp_var);
      add43_579 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_603_inst
    process(shl50_592, conv52_599) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_592, conv52_599, tmp_var);
      add53_604 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_628_inst
    process(shl60_617, conv62_624) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_617, conv62_624, tmp_var);
      add63_629 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_653_inst
    process(shl70_642, conv72_649) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_642, conv72_649, tmp_var);
      add73_654 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_478_inst
    process(shl_467, conv3_474) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_467, conv3_474, tmp_var);
      add_479 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1035_inst
    process(conv5x_xi_1031, elementx_x021x_xi_1005) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1031, elementx_x021x_xi_1005, tmp_var);
      addx_xi_1036 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1270_inst
    process(shl167_1259, conv170_1266) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1259, conv170_1266, tmp_var);
      add171_1271 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1288_inst
    process(shl173_1277, conv176_1284) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1277, conv176_1284, tmp_var);
      add177_1289 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1306_inst
    process(shl179_1295, conv182_1302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1295, conv182_1302, tmp_var);
      add183_1307 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1324_inst
    process(shl185_1313, conv188_1320) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1313, conv188_1320, tmp_var);
      add189_1325 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1342_inst
    process(shl191_1331, conv194_1338) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1331, conv194_1338, tmp_var);
      add195_1343 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1360_inst
    process(shl197_1349, conv200_1356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1349, conv200_1356, tmp_var);
      add201_1361 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1378_inst
    process(shl203_1367, conv206_1374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1367, conv206_1374, tmp_var);
      add207_1379 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1508_inst
    process(conv5x_xi364_1504, elementx_x021x_xi362_1478) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi364_1504, elementx_x021x_xi362_1478, tmp_var);
      addx_xi365_1509 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_801_inst
    process(shl92_790, conv95_797) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_790, conv95_797, tmp_var);
      add96_802 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_819_inst
    process(shl98_808, conv101_815) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_808, conv101_815, tmp_var);
      add102_820 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_837_inst
    process(shl104_826, conv107_833) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_826, conv107_833, tmp_var);
      add108_838 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_855_inst
    process(shl110_844, conv113_851) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_844, conv113_851, tmp_var);
      add114_856 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_873_inst
    process(shl116_862, conv119_869) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_862, conv119_869, tmp_var);
      add120_874 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_891_inst
    process(shl122_880, conv125_887) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_880, conv125_887, tmp_var);
      add126_892 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_909_inst
    process(shl128_898, conv131_905) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_898, conv131_905, tmp_var);
      add132_910 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_491_inst
    process(conv9_486) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_486, type_cast_490_wire_constant, tmp_var);
      shl10_492 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_516_inst
    process(conv19_511) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_511, type_cast_515_wire_constant, tmp_var);
      shl20_517 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_541_inst
    process(conv29_536) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_536, type_cast_540_wire_constant, tmp_var);
      shl30_542 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_566_inst
    process(conv39_561) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_561, type_cast_565_wire_constant, tmp_var);
      shl40_567 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_591_inst
    process(conv49_586) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_586, type_cast_590_wire_constant, tmp_var);
      shl50_592 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_616_inst
    process(conv59_611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_611, type_cast_615_wire_constant, tmp_var);
      shl60_617 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_641_inst
    process(conv69_636) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_636, type_cast_640_wire_constant, tmp_var);
      shl70_642 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_466_inst
    process(conv1_461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_461, type_cast_465_wire_constant, tmp_var);
      shl_467 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_988_inst
    process(mul82_672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_672, type_cast_987_wire_constant, tmp_var);
      conv2x_xi_989 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1041_inst
    process(addx_xi_1036) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1036, type_cast_1040_wire_constant, tmp_var);
      shl8x_xi_1042 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1068_inst
    process(conv83_678) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_678, type_cast_1067_wire_constant, tmp_var);
      Bx_xnot_1069 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1085_inst
    process(shl8x_xix_xlcssa_1059, sh_promx_xi_1081) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1059, sh_promx_xi_1081, tmp_var);
      shl14x_xi_1086 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1135_inst
    process(mul154_1130) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1130, type_cast_1134_wire_constant, tmp_var);
      sext_1136 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1258_inst
    process(conv165_1253) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1253, type_cast_1257_wire_constant, tmp_var);
      shl167_1259 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1276_inst
    process(add171_1271) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1271, type_cast_1275_wire_constant, tmp_var);
      shl173_1277 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1294_inst
    process(add177_1289) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1289, type_cast_1293_wire_constant, tmp_var);
      shl179_1295 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1312_inst
    process(add183_1307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1307, type_cast_1311_wire_constant, tmp_var);
      shl185_1313 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1330_inst
    process(add189_1325) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1325, type_cast_1329_wire_constant, tmp_var);
      shl191_1331 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1348_inst
    process(add195_1343) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1343, type_cast_1347_wire_constant, tmp_var);
      shl197_1349 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1366_inst
    process(add201_1361) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1361, type_cast_1365_wire_constant, tmp_var);
      shl203_1367 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1413_inst
    process(umax_1408) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1408, type_cast_1412_wire_constant, tmp_var);
      tmp414_1414 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1457_inst
    process(mul154_1130) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1130, type_cast_1456_wire_constant, tmp_var);
      iNsTr_55_1458 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1514_inst
    process(addx_xi365_1509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi365_1509, type_cast_1513_wire_constant, tmp_var);
      shl8x_xi366_1515 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1541_inst
    process(mul154_1130) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1130, type_cast_1540_wire_constant, tmp_var);
      iNsTr_87_1542 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1558_inst
    process(shl8x_xi366x_xlcssa_1532, sh_promx_xi375_1554) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi366x_xlcssa_1532, sh_promx_xi375_1554, tmp_var);
      shl14x_xi376_1559 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_789_inst
    process(conv90_784) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_784, type_cast_788_wire_constant, tmp_var);
      shl92_790 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_807_inst
    process(add96_802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_802, type_cast_806_wire_constant, tmp_var);
      shl98_808 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_825_inst
    process(add102_820) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_820, type_cast_824_wire_constant, tmp_var);
      shl104_826 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_843_inst
    process(add108_838) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_838, type_cast_842_wire_constant, tmp_var);
      shl110_844 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_861_inst
    process(add114_856) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_856, type_cast_860_wire_constant, tmp_var);
      shl116_862 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_879_inst
    process(add120_874) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_874, type_cast_878_wire_constant, tmp_var);
      shl122_880 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_897_inst
    process(add126_892) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_892, type_cast_896_wire_constant, tmp_var);
      shl128_898 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_944_inst
    process(umax427_939) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax427_939, type_cast_943_wire_constant, tmp_var);
      tmp428_945 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1727_inst
    process(conv289_1723, conv230_1715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv289_1723, conv230_1715, tmp_var);
      sub293_1728 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_683_inst
    process(mul82_672) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_672, type_cast_682_wire_constant, tmp_var);
      cmp387_684 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1150_inst
    process(conv155_1145) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1145, type_cast_1149_wire_constant, tmp_var);
      cmp161383_1151 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1169_inst
    process(tmp412_1164) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp412_1164, type_cast_1168_wire_constant, tmp_var);
      tmp413_1170 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1221_inst
    process(tmp22_1216) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp22_1216, type_cast_1220_wire_constant, tmp_var);
      tmp23_1222 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_717_inst
    process(tmp425_712) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp425_712, type_cast_716_wire_constant, tmp_var);
      tmp426_718 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_752_inst
    process(tmp30_747) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp30_747, type_cast_751_wire_constant, tmp_var);
      tmp31_753 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1050_inst
    process(convx_xi_1046, shlx_xi_995) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1046, shlx_xi_995, tmp_var);
      cmpx_xi_1051 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1523_inst
    process(convx_xi367_1519, shlx_xi359_1468) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi367_1519, shlx_xi359_1468, tmp_var);
      cmpx_xi368_1524 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1080_inst
    process(add1216x_xi_1075) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1075, type_cast_1079_wire_constant, tmp_var);
      sh_promx_xi_1081 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1553_inst
    process(add1216x_xi374_1548) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi374_1548, type_cast_1552_wire_constant, tmp_var);
      sh_promx_xi375_1554 <= tmp_var; --
    end process;
    -- shared split operator group (123) : array_obj_ref_1091_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1090_scaled;
      array_obj_ref_1091_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1091_index_offset_req_0;
      array_obj_ref_1091_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1091_index_offset_req_1;
      array_obj_ref_1091_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_1244_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar417_1243_scaled;
      array_obj_ref_1244_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1244_index_offset_req_0;
      array_obj_ref_1244_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1244_index_offset_req_1;
      array_obj_ref_1244_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_1564_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1563_scaled;
      array_obj_ref_1564_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1564_index_offset_req_0;
      array_obj_ref_1564_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1564_index_offset_req_1;
      array_obj_ref_1564_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- shared split operator group (126) : array_obj_ref_775_index_offset 
    ApIntAdd_group_126: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar431_774_scaled;
      array_obj_ref_775_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_775_index_offset_req_0;
      array_obj_ref_775_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_775_index_offset_req_1;
      array_obj_ref_775_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_126_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_126_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_126",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 126
    -- unary operator type_cast_1208_inst
    process(tmp20_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp20_1205, tmp_var);
      type_cast_1208_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1713_inst
    process(call229_1575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1575, tmp_var);
      type_cast_1713_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1721_inst
    process(call288_1718) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call288_1718, tmp_var);
      type_cast_1721_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_676_inst
    process(mul82_672) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_672, tmp_var);
      type_cast_676_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_704_inst
    process(tmp423_701) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp423_701, tmp_var);
      type_cast_704_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_739_inst
    process(tmp28_736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp28_736, tmp_var);
      type_cast_739_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1095_store_0 ptr_deref_912_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1095_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_912_store_0_req_0;
      ptr_deref_1095_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_912_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1095_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_912_store_0_req_1;
      ptr_deref_1095_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_912_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1095_word_address_0 & ptr_deref_912_word_address_0;
      data_in <= ptr_deref_1095_data_0 & ptr_deref_912_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1568_store_0 ptr_deref_1381_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1568_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1381_store_0_req_0;
      ptr_deref_1568_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1381_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1568_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1381_store_0_req_1;
      ptr_deref_1568_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1381_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1568_word_address_0 & ptr_deref_1381_word_address_0;
      data_in <= ptr_deref_1568_data_0 & ptr_deref_1381_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_456_inst RPIPE_maxpool_input_pipe_544_inst RPIPE_maxpool_input_pipe_606_inst RPIPE_maxpool_input_pipe_581_inst RPIPE_maxpool_input_pipe_494_inst RPIPE_maxpool_input_pipe_556_inst RPIPE_maxpool_input_pipe_631_inst RPIPE_maxpool_input_pipe_519_inst RPIPE_maxpool_input_pipe_619_inst RPIPE_maxpool_input_pipe_469_inst RPIPE_maxpool_input_pipe_481_inst RPIPE_maxpool_input_pipe_569_inst RPIPE_maxpool_input_pipe_644_inst RPIPE_maxpool_input_pipe_506_inst RPIPE_maxpool_input_pipe_594_inst RPIPE_maxpool_input_pipe_531_inst RPIPE_maxpool_input_pipe_1297_inst RPIPE_maxpool_input_pipe_1333_inst RPIPE_maxpool_input_pipe_1279_inst RPIPE_maxpool_input_pipe_1248_inst RPIPE_maxpool_input_pipe_1261_inst RPIPE_maxpool_input_pipe_1351_inst RPIPE_maxpool_input_pipe_1369_inst RPIPE_maxpool_input_pipe_1315_inst RPIPE_maxpool_input_pipe_1499_inst RPIPE_maxpool_input_pipe_779_inst RPIPE_maxpool_input_pipe_792_inst RPIPE_maxpool_input_pipe_810_inst RPIPE_maxpool_input_pipe_828_inst RPIPE_maxpool_input_pipe_846_inst RPIPE_maxpool_input_pipe_864_inst RPIPE_maxpool_input_pipe_882_inst RPIPE_maxpool_input_pipe_900_inst RPIPE_maxpool_input_pipe_1026_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_456_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_544_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_606_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_581_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_494_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_556_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_631_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_519_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_619_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_469_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_481_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_569_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_644_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_506_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_594_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_531_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1297_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1333_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1279_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1248_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1261_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_1351_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1369_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1315_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1499_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_779_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_792_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_810_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_828_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_846_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_864_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_882_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_900_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1026_inst_req_0;
      RPIPE_maxpool_input_pipe_456_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_544_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_606_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_581_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_494_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_556_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_631_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_519_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_619_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_469_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_481_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_569_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_644_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_506_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_594_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_531_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1297_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1333_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1279_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1248_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1261_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_1351_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1369_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1315_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1499_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_779_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_792_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_810_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_828_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_846_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_864_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_882_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_900_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1026_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_456_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_544_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_606_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_581_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_494_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_556_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_631_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_519_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_619_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_469_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_481_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_569_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_644_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_506_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_594_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_531_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1297_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1333_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1279_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1248_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1261_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_1351_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1369_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1315_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1499_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_779_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_792_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_810_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_828_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_846_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_864_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_882_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_900_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1026_inst_req_1;
      RPIPE_maxpool_input_pipe_456_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_544_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_606_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_581_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_494_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_556_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_631_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_519_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_619_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_469_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_481_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_569_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_644_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_506_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_594_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_531_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1297_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1333_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1279_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1248_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1261_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_1351_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1369_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1315_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1499_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_779_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_792_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_810_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_828_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_846_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_864_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_882_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_900_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1026_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call_457 <= data_out(271 downto 264);
      call31_545 <= data_out(263 downto 256);
      call56_607 <= data_out(255 downto 248);
      call46_582 <= data_out(247 downto 240);
      call11_495 <= data_out(239 downto 232);
      call36_557 <= data_out(231 downto 224);
      call66_632 <= data_out(223 downto 216);
      call21_520 <= data_out(215 downto 208);
      call61_620 <= data_out(207 downto 200);
      call2_470 <= data_out(199 downto 192);
      call6_482 <= data_out(191 downto 184);
      call41_570 <= data_out(183 downto 176);
      call71_645 <= data_out(175 downto 168);
      call16_507 <= data_out(167 downto 160);
      call51_595 <= data_out(159 downto 152);
      call26_532 <= data_out(151 downto 144);
      call180_1298 <= data_out(143 downto 136);
      call192_1334 <= data_out(135 downto 128);
      call174_1280 <= data_out(127 downto 120);
      call164_1249 <= data_out(119 downto 112);
      call168_1262 <= data_out(111 downto 104);
      call198_1352 <= data_out(103 downto 96);
      call204_1370 <= data_out(95 downto 88);
      call186_1316 <= data_out(87 downto 80);
      callx_xi363_1500 <= data_out(79 downto 72);
      call89_780 <= data_out(71 downto 64);
      call93_793 <= data_out(63 downto 56);
      call99_811 <= data_out(55 downto 48);
      call105_829 <= data_out(47 downto 40);
      call111_847 <= data_out(39 downto 32);
      call117_865 <= data_out(31 downto 24);
      call123_883 <= data_out(23 downto 16);
      call129_901 <= data_out(15 downto 8);
      callx_xi_1027 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1582_inst WPIPE_maxpool_output_pipe_1586_inst WPIPE_maxpool_output_pipe_1818_inst WPIPE_maxpool_output_pipe_1803_inst WPIPE_maxpool_output_pipe_1806_inst WPIPE_maxpool_output_pipe_1812_inst WPIPE_maxpool_output_pipe_1821_inst WPIPE_maxpool_output_pipe_1809_inst WPIPE_maxpool_output_pipe_1815_inst WPIPE_maxpool_output_pipe_1824_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1582_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1586_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1818_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1803_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1806_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1812_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1821_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1809_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1815_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1824_inst_req_0;
      WPIPE_maxpool_output_pipe_1582_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1586_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1818_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1803_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1806_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1812_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1821_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1809_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1815_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1824_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1582_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1586_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1818_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1803_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1806_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1812_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1821_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1809_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1815_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1824_inst_req_1;
      WPIPE_maxpool_output_pipe_1582_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1586_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1818_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1803_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1806_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1812_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1821_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1809_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1815_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1824_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= type_cast_1584_wire_constant & type_cast_1588_wire_constant & conv309_1752 & conv339_1802 & conv333_1792 & conv321_1772 & conv303_1742 & conv327_1782 & conv315_1762 & conv297_1732;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_1665_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1665_inst_req_0;
      WPIPE_num_out_pipe_1665_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1665_inst_req_1;
      WPIPE_num_out_pipe_1665_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul249_1594;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1575_call call_stmt_1718_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1575_call_req_0;
      reqL_unguarded(0) <= call_stmt_1718_call_req_0;
      call_stmt_1575_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1718_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1575_call_req_1;
      reqR_unguarded(0) <= call_stmt_1718_call_req_1;
      call_stmt_1575_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1718_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_1575 <= data_out(127 downto 64);
      call288_1718 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1685_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(135 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1685_call_req_0;
      call_stmt_1685_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1685_call_req_1;
      call_stmt_1685_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv255_1671 & conv261_1675 & and264_1681;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 136,
        owidth => 136,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(135 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1692_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1692_call_req_0;
      call_stmt_1692_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1692_call_req_1;
      call_stmt_1692_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul236_1581 & add33_554 & sub_1600 & sub273_1606 & add23_529 & add13_504;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4061_start: Boolean;
  signal convolve_CP_4061_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_input_done_pipe_1982_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1875_inst_req_1 : boolean;
  signal type_cast_1999_inst_req_0 : boolean;
  signal slice_1991_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1997_inst_req_1 : boolean;
  signal NOT_u1_u1_1942_inst_ack_0 : boolean;
  signal W_next_sum_1971_delayed_1_0_2001_inst_req_0 : boolean;
  signal NOT_u1_u1_1942_inst_req_0 : boolean;
  signal type_cast_1999_inst_ack_0 : boolean;
  signal type_cast_2007_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1875_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2005_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_1887_inst_ack_0 : boolean;
  signal n_out_count_1975_1870_buf_req_0 : boolean;
  signal RPIPE_kernel_pipe2_1887_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2005_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1875_inst_req_0 : boolean;
  signal phi_stmt_1868_req_1 : boolean;
  signal SUB_u31_u31_1907_inst_ack_1 : boolean;
  signal type_cast_2007_inst_ack_0 : boolean;
  signal phi_stmt_1868_ack_0 : boolean;
  signal slice_1991_inst_ack_0 : boolean;
  signal n_out_count_1975_1870_buf_ack_0 : boolean;
  signal nacc_1926_1867_buf_req_0 : boolean;
  signal W_next_sum_1971_delayed_1_0_2001_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1997_inst_ack_1 : boolean;
  signal slice_1991_inst_req_1 : boolean;
  signal NOT_u1_u1_1942_inst_req_1 : boolean;
  signal nacc_1926_1867_buf_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2005_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1875_inst_ack_1 : boolean;
  signal slice_1991_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1997_inst_ack_0 : boolean;
  signal type_cast_2007_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_1887_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1883_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1883_inst_ack_0 : boolean;
  signal n_out_count_1975_1870_buf_req_1 : boolean;
  signal W_next_sum_1971_delayed_1_0_2001_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_1887_inst_ack_1 : boolean;
  signal NOT_u1_u1_1942_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2005_inst_ack_0 : boolean;
  signal n_out_count_1975_1870_buf_ack_1 : boolean;
  signal type_cast_1999_inst_req_1 : boolean;
  signal type_cast_2007_inst_ack_1 : boolean;
  signal slice_1987_inst_req_0 : boolean;
  signal W_next_sum_1971_delayed_1_0_2001_inst_ack_1 : boolean;
  signal type_cast_1999_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1883_inst_req_1 : boolean;
  signal W_next_sum_1966_delayed_1_0_1993_inst_req_0 : boolean;
  signal do_while_stmt_1858_branch_ack_0 : boolean;
  signal W_next_sum_1966_delayed_1_0_1993_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1883_inst_ack_1 : boolean;
  signal W_next_sum_1966_delayed_1_0_1993_inst_req_1 : boolean;
  signal W_next_sum_1966_delayed_1_0_1993_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1997_inst_req_0 : boolean;
  signal SUB_u31_u31_1907_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1957_inst_req_0 : boolean;
  signal SUB_u31_u31_1907_inst_ack_0 : boolean;
  signal nacc_1926_1867_buf_req_1 : boolean;
  signal nacc_1926_1867_buf_ack_1 : boolean;
  signal do_while_stmt_1858_branch_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1957_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_1961_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_1961_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe2_1961_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_1961_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1957_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1957_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1836_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1836_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1836_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1836_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1839_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1839_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1839_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1839_inst_ack_1 : boolean;
  signal slice_1843_inst_req_0 : boolean;
  signal slice_1843_inst_ack_0 : boolean;
  signal slice_1843_inst_req_1 : boolean;
  signal slice_1843_inst_ack_1 : boolean;
  signal slice_1847_inst_req_0 : boolean;
  signal slice_1847_inst_ack_0 : boolean;
  signal slice_1847_inst_req_1 : boolean;
  signal slice_1847_inst_ack_1 : boolean;
  signal SUB_u31_u31_1907_inst_req_1 : boolean;
  signal phi_stmt_1868_req_0 : boolean;
  signal WPIPE_input_done_pipe_1982_inst_req_1 : boolean;
  signal do_while_stmt_1858_branch_req_0 : boolean;
  signal WPIPE_input_done_pipe_1982_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_1982_inst_req_0 : boolean;
  signal phi_stmt_1860_req_1 : boolean;
  signal slice_1987_inst_ack_1 : boolean;
  signal slice_1987_inst_req_1 : boolean;
  signal phi_stmt_1860_req_0 : boolean;
  signal phi_stmt_1860_ack_0 : boolean;
  signal slice_1987_inst_ack_0 : boolean;
  signal nmycount_1934_1863_buf_req_0 : boolean;
  signal nmycount_1934_1863_buf_ack_0 : boolean;
  signal nmycount_1934_1863_buf_req_1 : boolean;
  signal nmycount_1934_1863_buf_ack_1 : boolean;
  signal phi_stmt_1864_req_1 : boolean;
  signal phi_stmt_1864_req_0 : boolean;
  signal phi_stmt_1864_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4061_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4061_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4061_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4061_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4061: Block -- control-path 
    signal convolve_CP_4061_elements: BooleanArray(144 downto 0);
    -- 
  begin -- 
    convolve_CP_4061_elements(0) <= convolve_CP_4061_start;
    convolve_CP_4061_symbol <= convolve_CP_4061_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	144 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1833/merge_stmt_1834_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1833/merge_stmt_1834__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1833/merge_stmt_1834__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_1833/$entry
      -- CP-element group 0: 	 branch_block_stmt_1833/branch_block_stmt_1833__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1833/merge_stmt_1834__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1833/branch_block_stmt_1833__exit__
      -- CP-element group 1: 	 branch_block_stmt_1833/$exit
      -- CP-element group 1: 	 $exit
      -- 
    convolve_CP_4061_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	143 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	144 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1833/do_while_stmt_1858__exit__
      -- CP-element group 2: 	 branch_block_stmt_1833/loopback
      -- CP-element group 2: 	 branch_block_stmt_1833/loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1833/loopback_PhiReq/$exit
      -- 
    convolve_CP_4061_elements(2) <= convolve_CP_4061_elements(143);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	144 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Update/cr
      -- 
    ra_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1836_inst_ack_0, ack => convolve_CP_4061_elements(3)); -- 
    cr_4091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(3), ack => RPIPE_num_out_pipe_1836_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Update/ca
      -- 
    ca_4092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1836_inst_ack_1, ack => convolve_CP_4061_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	144 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Update/cr
      -- 
    ra_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1839_inst_ack_0, ack => convolve_CP_4061_elements(5)); -- 
    cr_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(5), ack => RPIPE_size_pipe_1839_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Sample/rr
      -- 
    ca_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1839_inst_ack_1, ack => convolve_CP_4061_elements(6)); -- 
    rr_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(6), ack => slice_1847_inst_req_0); -- 
    rr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(6), ack => slice_1843_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Sample/ra
      -- 
    ra_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1843_inst_ack_0, ack => convolve_CP_4061_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	144 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Update/ca
      -- 
    ca_4120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1843_inst_ack_1, ack => convolve_CP_4061_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Sample/ra
      -- 
    ra_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1847_inst_ack_0, ack => convolve_CP_4061_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	144 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Update/ca
      -- 
    ca_4134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1847_inst_ack_1, ack => convolve_CP_4061_elements(10)); -- 
    -- CP-element group 11:  join  transition  place  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	4 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/$exit
      -- CP-element group 11: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857__exit__
      -- CP-element group 11: 	 branch_block_stmt_1833/do_while_stmt_1858__entry__
      -- 
    convolve_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(10) & convolve_CP_4061_elements(8) & convolve_CP_4061_elements(4);
      gj_convolve_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	18 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1833/do_while_stmt_1858/$entry
      -- CP-element group 12: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858__entry__
      -- 
    convolve_CP_4061_elements(12) <= convolve_CP_4061_elements(11);
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	143 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858__exit__
      -- 
    -- Element group convolve_CP_4061_elements(13) is bound as output of CP function.
    -- CP-element group 14:  merge  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_back
      -- 
    -- Element group convolve_CP_4061_elements(14) is bound as output of CP function.
    -- CP-element group 15:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	141 
    -- CP-element group 15: 	142 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_exit/$entry
      -- CP-element group 15: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_taken/$entry
      -- CP-element group 15: 	 branch_block_stmt_1833/do_while_stmt_1858/condition_done
      -- 
    convolve_CP_4061_elements(15) <= convolve_CP_4061_elements(20);
    -- CP-element group 16:  branch  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	140 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_body_done
      -- 
    convolve_CP_4061_elements(16) <= convolve_CP_4061_elements(140);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	67 
    -- CP-element group 17: 	50 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4061_elements(17) <= convolve_CP_4061_elements(14);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	69 
    -- CP-element group 18: 	52 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4061_elements(18) <= convolve_CP_4061_elements(12);
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	64 
    -- CP-element group 19: 	25 
    -- CP-element group 19: 	26 
    -- CP-element group 19: 	139 
    -- CP-element group 19: 	88 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	45 
    -- CP-element group 19: 	92 
    -- CP-element group 19: 	96 
    -- CP-element group 19: 	80 
    -- CP-element group 19: 	84 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/$entry
      -- CP-element group 19: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_4061_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	66 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	139 
    -- CP-element group 20: 	30 
    -- CP-element group 20: 	95 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/condition_evaluated
      -- 
    condition_evaluated_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(20), ack => do_while_stmt_1858_branch_req_0); -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(66) & convolve_CP_4061_elements(24) & convolve_CP_4061_elements(139) & convolve_CP_4061_elements(30) & convolve_CP_4061_elements(95);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	63 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	44 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	46 
    -- CP-element group 21: 	27 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(63) & convolve_CP_4061_elements(25) & convolve_CP_4061_elements(44) & convolve_CP_4061_elements(24);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	65 
    -- CP-element group 22: 	47 
    -- CP-element group 22: 	28 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	85 
    -- CP-element group 22: 	89 
    -- CP-element group 22: 	93 
    -- CP-element group 22: 	81 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	63 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	44 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/aggregated_phi_sample_ack
      -- CP-element group 22: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_sample_completed_
      -- 
    convolve_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(65) & convolve_CP_4061_elements(47) & convolve_CP_4061_elements(28);
      gj_convolve_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	64 
    -- CP-element group 23: 	26 
    -- CP-element group 23: 	45 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23: 	29 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/aggregated_phi_update_req
      -- CP-element group 23: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_update_start__ps
      -- 
    convolve_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(64) & convolve_CP_4061_elements(26) & convolve_CP_4061_elements(45);
      gj_convolve_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	66 
    -- CP-element group 24: 	49 
    -- CP-element group 24: 	30 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	21 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(66) & convolve_CP_4061_elements(49) & convolve_CP_4061_elements(30);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	19 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: 	95 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	21 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_sample_start_
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(22) & convolve_CP_4061_elements(95);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	130 
    -- CP-element group 26: 	119 
    -- CP-element group 26: 	30 
    -- CP-element group 26: 	107 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	23 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_update_start_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(130) & convolve_CP_4061_elements(119) & convolve_CP_4061_elements(30) & convolve_CP_4061_elements(107);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	21 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_sample_start__ps
      -- 
    convolve_CP_4061_elements(27) <= convolve_CP_4061_elements(21);
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	22 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_sample_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_update_start__ps
      -- 
    convolve_CP_4061_elements(29) <= convolve_CP_4061_elements(23);
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: 	128 
    -- CP-element group 30: 	117 
    -- CP-element group 30: 	20 
    -- CP-element group 30: 	106 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	26 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_update_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	17 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_loopback_trigger
      -- 
    convolve_CP_4061_elements(31) <= convolve_CP_4061_elements(17);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_loopback_sample_req
      -- CP-element group 32: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_loopback_sample_req_ps
      -- 
    phi_stmt_1860_loopback_sample_req_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_loopback_sample_req_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(32), ack => phi_stmt_1860_req_1); -- 
    -- Element group convolve_CP_4061_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	18 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_entry_trigger
      -- 
    convolve_CP_4061_elements(33) <= convolve_CP_4061_elements(18);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_entry_sample_req
      -- CP-element group 34: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_entry_sample_req_ps
      -- 
    phi_stmt_1860_entry_sample_req_4167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_entry_sample_req_4167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(34), ack => phi_stmt_1860_req_0); -- 
    -- Element group convolve_CP_4061_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_phi_mux_ack
      -- CP-element group 35: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1860_phi_mux_ack_ps
      -- 
    phi_stmt_1860_phi_mux_ack_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1860_ack_0, ack => convolve_CP_4061_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_sample_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_sample_completed_
      -- 
    -- Element group convolve_CP_4061_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_update_start__ps
      -- CP-element group 37: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_update_start_
      -- 
    -- Element group convolve_CP_4061_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_update_completed__ps
      -- 
    convolve_CP_4061_elements(38) <= convolve_CP_4061_elements(39);
    -- CP-element group 39:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	38 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_mcount_var_1862_update_completed_
      -- 
    -- Element group convolve_CP_4061_elements(39) is a control-delay.
    cp_element_39_delay: control_delay_element  generic map(name => " 39_delay", delay_value => 1)  port map(req => convolve_CP_4061_elements(37), ack => convolve_CP_4061_elements(39), clk => clk, reset =>reset);
    -- CP-element group 40:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_sample_start__ps
      -- CP-element group 40: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Sample/req
      -- 
    req_4191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(40), ack => nmycount_1934_1863_buf_req_0); -- 
    -- Element group convolve_CP_4061_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_update_start__ps
      -- CP-element group 41: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Update/req
      -- 
    req_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(41), ack => nmycount_1934_1863_buf_req_1); -- 
    -- Element group convolve_CP_4061_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_sample_completed__ps
      -- CP-element group 42: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Sample/ack
      -- 
    ack_4192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1934_1863_buf_ack_0, ack => convolve_CP_4061_elements(42)); -- 
    -- CP-element group 43:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_update_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nmycount_1863_Update/ack
      -- 
    ack_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1934_1863_buf_ack_1, ack => convolve_CP_4061_elements(43)); -- 
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	22 
    -- CP-element group 44: 	87 
    -- CP-element group 44: 	91 
    -- CP-element group 44: 	95 
    -- CP-element group 44: 	83 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_sample_start_
      -- 
    convolve_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(22) & convolve_CP_4061_elements(87) & convolve_CP_4061_elements(91) & convolve_CP_4061_elements(95) & convolve_CP_4061_elements(83);
      gj_convolve_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	19 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	111 
    -- CP-element group 45: 	115 
    -- CP-element group 45: 	49 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	23 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_update_start_
      -- 
    convolve_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(111) & convolve_CP_4061_elements(115) & convolve_CP_4061_elements(49);
      gj_convolve_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	21 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_sample_start__ps
      -- 
    convolve_CP_4061_elements(46) <= convolve_CP_4061_elements(21);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	22 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_sample_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(47) is bound as output of CP function.
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_update_start__ps
      -- 
    convolve_CP_4061_elements(48) <= convolve_CP_4061_elements(23);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	24 
    -- CP-element group 49: 	109 
    -- CP-element group 49: 	113 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	45 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_update_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	17 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_loopback_trigger
      -- 
    convolve_CP_4061_elements(50) <= convolve_CP_4061_elements(17);
    -- CP-element group 51:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_loopback_sample_req
      -- CP-element group 51: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_loopback_sample_req_ps
      -- 
    phi_stmt_1864_loopback_sample_req_4208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1864_loopback_sample_req_4208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(51), ack => phi_stmt_1864_req_1); -- 
    -- Element group convolve_CP_4061_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	18 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_entry_trigger
      -- 
    convolve_CP_4061_elements(52) <= convolve_CP_4061_elements(18);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_entry_sample_req
      -- CP-element group 53: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_entry_sample_req_ps
      -- 
    phi_stmt_1864_entry_sample_req_4211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1864_entry_sample_req_4211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(53), ack => phi_stmt_1864_req_0); -- 
    -- Element group convolve_CP_4061_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_phi_mux_ack
      -- CP-element group 54: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1864_phi_mux_ack_ps
      -- 
    phi_stmt_1864_phi_mux_ack_4214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1864_ack_0, ack => convolve_CP_4061_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_sample_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_update_start__ps
      -- 
    -- Element group convolve_CP_4061_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_update_completed__ps
      -- 
    convolve_CP_4061_elements(57) <= convolve_CP_4061_elements(58);
    -- CP-element group 58:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	57 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_acc_var_1866_update_completed_
      -- 
    -- Element group convolve_CP_4061_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => convolve_CP_4061_elements(56), ack => convolve_CP_4061_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Sample/req
      -- 
    req_4235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(59), ack => nacc_1926_1867_buf_req_0); -- 
    -- Element group convolve_CP_4061_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_update_start__ps
      -- CP-element group 60: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Update/req
      -- 
    req_4240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(60), ack => nacc_1926_1867_buf_req_1); -- 
    -- Element group convolve_CP_4061_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_sample_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Sample/ack
      -- 
    ack_4236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1926_1867_buf_ack_0, ack => convolve_CP_4061_elements(61)); -- 
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_nacc_1867_Update/ack
      -- 
    ack_4241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1926_1867_buf_ack_1, ack => convolve_CP_4061_elements(62)); -- 
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	22 
    -- CP-element group 63: 	95 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	21 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_sample_start_
      -- 
    convolve_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(22) & convolve_CP_4061_elements(95);
      gj_convolve_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	19 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	101 
    -- CP-element group 64: 	104 
    -- CP-element group 64: 	107 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	23 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_update_start_
      -- 
    convolve_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(66) & convolve_CP_4061_elements(101) & convolve_CP_4061_elements(104) & convolve_CP_4061_elements(107);
      gj_convolve_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	22 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_sample_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	24 
    -- CP-element group 66: 	20 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	106 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_update_completed__ps
      -- 
    -- Element group convolve_CP_4061_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	17 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_loopback_trigger
      -- 
    convolve_CP_4061_elements(67) <= convolve_CP_4061_elements(17);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_loopback_sample_req_ps
      -- CP-element group 68: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_loopback_sample_req
      -- 
    phi_stmt_1868_loopback_sample_req_4252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_loopback_sample_req_4252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(68), ack => phi_stmt_1868_req_0); -- 
    -- Element group convolve_CP_4061_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	18 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_entry_trigger
      -- 
    convolve_CP_4061_elements(69) <= convolve_CP_4061_elements(18);
    -- CP-element group 70:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_entry_sample_req_ps
      -- CP-element group 70: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_entry_sample_req
      -- 
    phi_stmt_1868_entry_sample_req_4255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1868_entry_sample_req_4255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(70), ack => phi_stmt_1868_req_1); -- 
    -- Element group convolve_CP_4061_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_phi_mux_ack
      -- CP-element group 71: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/phi_stmt_1868_phi_mux_ack_ps
      -- 
    phi_stmt_1868_phi_mux_ack_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1868_ack_0, ack => convolve_CP_4061_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Sample/req
      -- CP-element group 72: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_sample_start_
      -- 
    req_4271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(72), ack => n_out_count_1975_1870_buf_req_0); -- 
    -- Element group convolve_CP_4061_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Update/req
      -- CP-element group 73: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_update_start__ps
      -- 
    req_4276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(73), ack => n_out_count_1975_1870_buf_req_1); -- 
    -- Element group convolve_CP_4061_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Sample/ack
      -- CP-element group 74: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_sample_completed__ps
      -- 
    ack_4272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1975_1870_buf_ack_0, ack => convolve_CP_4061_elements(74)); -- 
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_Update/ack
      -- CP-element group 75: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/R_n_out_count_1870_update_completed__ps
      -- 
    ack_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1975_1870_buf_ack_1, ack => convolve_CP_4061_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_sample_start__ps
      -- CP-element group 76: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_sample_start_
      -- 
    -- Element group convolve_CP_4061_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_update_start__ps
      -- 
    -- Element group convolve_CP_4061_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_update_completed__ps
      -- 
    convolve_CP_4061_elements(78) <= convolve_CP_4061_elements(79);
    -- CP-element group 79:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1872_update_completed_
      -- 
    -- Element group convolve_CP_4061_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convolve_CP_4061_elements(77), ack => convolve_CP_4061_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	19 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	83 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_sample_start_
      -- 
    rr_4294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(80), ack => RPIPE_input_pipe1_1875_inst_req_0); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(83);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	22 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	111 
    -- CP-element group 81: 	115 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_update_start_
      -- 
    cr_4299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(81), ack => RPIPE_input_pipe1_1875_inst_req_1); -- 
    convolve_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(22) & convolve_CP_4061_elements(82) & convolve_CP_4061_elements(111) & convolve_CP_4061_elements(115);
      gj_convolve_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	81 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_sample_completed_
      -- 
    ra_4295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1875_inst_ack_0, ack => convolve_CP_4061_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	109 
    -- CP-element group 83: 	113 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	44 
    -- CP-element group 83: 	80 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_input_pipe1_1875_update_completed_
      -- 
    ca_4300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1875_inst_ack_1, ack => convolve_CP_4061_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	19 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	87 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_sample_start_
      -- 
    rr_4308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(84), ack => RPIPE_kernel_pipe1_1883_inst_req_0); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(87);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	22 
    -- CP-element group 85: 	86 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	111 
    -- CP-element group 85: 	115 
    -- CP-element group 85: 	101 
    -- CP-element group 85: 	104 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Update/cr
      -- 
    cr_4313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(85), ack => RPIPE_kernel_pipe1_1883_inst_req_1); -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(22) & convolve_CP_4061_elements(86) & convolve_CP_4061_elements(111) & convolve_CP_4061_elements(115) & convolve_CP_4061_elements(101) & convolve_CP_4061_elements(104);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	85 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_sample_completed_
      -- 
    ra_4309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1883_inst_ack_0, ack => convolve_CP_4061_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	109 
    -- CP-element group 87: 	113 
    -- CP-element group 87: 	100 
    -- CP-element group 87: 	103 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	44 
    -- CP-element group 87: 	84 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe1_1883_Update/ca
      -- 
    ca_4314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1883_inst_ack_1, ack => convolve_CP_4061_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	19 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	91 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Sample/$entry
      -- 
    rr_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(88), ack => RPIPE_kernel_pipe2_1887_inst_req_0); -- 
    convolve_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(91);
      gj_convolve_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	22 
    -- CP-element group 89: 	90 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	111 
    -- CP-element group 89: 	115 
    -- CP-element group 89: 	101 
    -- CP-element group 89: 	104 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Update/cr
      -- CP-element group 89: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_update_start_
      -- 
    cr_4327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(89), ack => RPIPE_kernel_pipe2_1887_inst_req_1); -- 
    convolve_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(22) & convolve_CP_4061_elements(90) & convolve_CP_4061_elements(111) & convolve_CP_4061_elements(115) & convolve_CP_4061_elements(101) & convolve_CP_4061_elements(104);
      gj_convolve_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Sample/$exit
      -- 
    ra_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_1887_inst_ack_0, ack => convolve_CP_4061_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	109 
    -- CP-element group 91: 	113 
    -- CP-element group 91: 	100 
    -- CP-element group 91: 	103 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: 	44 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/RPIPE_kernel_pipe2_1887_update_completed_
      -- 
    ca_4328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_1887_inst_ack_1, ack => convolve_CP_4061_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	19 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Sample/rr
      -- 
    rr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(92), ack => SUB_u31_u31_1907_inst_req_0); -- 
    convolve_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(94);
      gj_convolve_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	22 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	130 
    -- CP-element group 93: 	119 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	107 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_update_start_
      -- CP-element group 93: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Update/cr
      -- 
    cr_4341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(93), ack => SUB_u31_u31_1907_inst_req_1); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(22) & convolve_CP_4061_elements(130) & convolve_CP_4061_elements(119) & convolve_CP_4061_elements(95) & convolve_CP_4061_elements(107);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Sample/ra
      -- 
    ra_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u31_u31_1907_inst_ack_0, ack => convolve_CP_4061_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	128 
    -- CP-element group 95: 	117 
    -- CP-element group 95: 	20 
    -- CP-element group 95: 	106 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	63 
    -- CP-element group 95: 	25 
    -- CP-element group 95: 	44 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/SUB_u31_u31_1907_Update/$exit
      -- 
    ca_4342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u31_u31_1907_inst_ack_1, ack => convolve_CP_4061_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	19 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Sample/rr
      -- 
    rr_4350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(96), ack => NOT_u1_u1_1942_inst_req_0); -- 
    convolve_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(19) & convolve_CP_4061_elements(98);
      gj_convolve_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	101 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_update_start_
      -- CP-element group 97: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Update/cr
      -- 
    cr_4355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(97), ack => NOT_u1_u1_1942_inst_req_1); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(99) & convolve_CP_4061_elements(101);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_sample_completed_
      -- 
    ra_4351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1942_inst_ack_0, ack => convolve_CP_4061_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/NOT_u1_u1_1942_update_completed_
      -- 
    ca_4356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1942_inst_ack_1, ack => convolve_CP_4061_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: 	87 
    -- CP-element group 100: 	91 
    -- CP-element group 100: 	99 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Sample/req
      -- 
    req_4364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(100), ack => WPIPE_kernel_pipe1_1957_inst_req_0); -- 
    convolve_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(66) & convolve_CP_4061_elements(87) & convolve_CP_4061_elements(91) & convolve_CP_4061_elements(99) & convolve_CP_4061_elements(102);
      gj_convolve_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	64 
    -- CP-element group 101: 	85 
    -- CP-element group 101: 	89 
    -- CP-element group 101: 	97 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Update/req
      -- CP-element group 101: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Update/$entry
      -- 
    ack_4365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1957_inst_ack_0, ack => convolve_CP_4061_elements(101)); -- 
    req_4369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(101), ack => WPIPE_kernel_pipe1_1957_inst_req_1); -- 
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	140 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe1_1957_Update/$exit
      -- 
    ack_4370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1957_inst_ack_1, ack => convolve_CP_4061_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: 	87 
    -- CP-element group 103: 	91 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Sample/req
      -- CP-element group 103: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_sample_start_
      -- 
    req_4378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(103), ack => WPIPE_kernel_pipe2_1961_inst_req_0); -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(66) & convolve_CP_4061_elements(87) & convolve_CP_4061_elements(91) & convolve_CP_4061_elements(105);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	64 
    -- CP-element group 104: 	85 
    -- CP-element group 104: 	89 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Sample/ack
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_sample_completed_
      -- 
    ack_4379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_1961_inst_ack_0, ack => convolve_CP_4061_elements(104)); -- 
    req_4383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(104), ack => WPIPE_kernel_pipe2_1961_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	140 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	103 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Update/ack
      -- CP-element group 105: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_kernel_pipe2_1961_update_completed_
      -- 
    ack_4384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_1961_inst_ack_1, ack => convolve_CP_4061_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: 	30 
    -- CP-element group 106: 	95 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Sample/req
      -- 
    req_4392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(106), ack => WPIPE_input_done_pipe_1982_inst_req_0); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(66) & convolve_CP_4061_elements(30) & convolve_CP_4061_elements(95) & convolve_CP_4061_elements(108);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	64 
    -- CP-element group 107: 	26 
    -- CP-element group 107: 	93 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Update/req
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Sample/ack
      -- 
    ack_4393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1982_inst_ack_0, ack => convolve_CP_4061_elements(107)); -- 
    req_4397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(107), ack => WPIPE_input_done_pipe_1982_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	140 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Update/ack
      -- CP-element group 108: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_input_done_pipe_1982_Update/$exit
      -- 
    ack_4398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1982_inst_ack_1, ack => convolve_CP_4061_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	87 
    -- CP-element group 109: 	49 
    -- CP-element group 109: 	91 
    -- CP-element group 109: 	83 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Sample/rr
      -- 
    rr_4406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(109), ack => slice_1987_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 15,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(87) & convolve_CP_4061_elements(49) & convolve_CP_4061_elements(91) & convolve_CP_4061_elements(83) & convolve_CP_4061_elements(111);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	123 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Update/cr
      -- 
    cr_4411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(110), ack => slice_1987_inst_req_1); -- 
    convolve_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(123) & convolve_CP_4061_elements(112);
      gj_convolve_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	85 
    -- CP-element group 111: 	89 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	45 
    -- CP-element group 111: 	81 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Sample/ra
      -- 
    ra_4407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1987_inst_ack_0, ack => convolve_CP_4061_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	121 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1987_Update/ca
      -- 
    ca_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1987_inst_ack_1, ack => convolve_CP_4061_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	87 
    -- CP-element group 113: 	49 
    -- CP-element group 113: 	91 
    -- CP-element group 113: 	83 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_sample_start_
      -- 
    rr_4420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(113), ack => slice_1991_inst_req_0); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 15,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(87) & convolve_CP_4061_elements(49) & convolve_CP_4061_elements(91) & convolve_CP_4061_elements(83) & convolve_CP_4061_elements(115);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	134 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_update_start_
      -- 
    cr_4425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(114), ack => slice_1991_inst_req_1); -- 
    convolve_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(134) & convolve_CP_4061_elements(116);
      gj_convolve_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	85 
    -- CP-element group 115: 	89 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	45 
    -- CP-element group 115: 	81 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_sample_completed_
      -- 
    ra_4421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1991_inst_ack_0, ack => convolve_CP_4061_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	132 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/slice_1991_update_completed_
      -- 
    ca_4426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1991_inst_ack_1, ack => convolve_CP_4061_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	30 
    -- CP-element group 117: 	95 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Sample/req
      -- 
    req_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(117), ack => W_next_sum_1966_delayed_1_0_1993_inst_req_0); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(30) & convolve_CP_4061_elements(95) & convolve_CP_4061_elements(119);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	123 
    -- CP-element group 118: 	126 
    -- CP-element group 118: 	120 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_update_start_
      -- CP-element group 118: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Update/req
      -- 
    req_4439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(118), ack => W_next_sum_1966_delayed_1_0_1993_inst_req_1); -- 
    convolve_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(123) & convolve_CP_4061_elements(126) & convolve_CP_4061_elements(120);
      gj_convolve_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	26 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	93 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Sample/ack
      -- 
    ack_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1966_delayed_1_0_1993_inst_ack_0, ack => convolve_CP_4061_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	125 
    -- CP-element group 120: 	121 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_1995_Update/ack
      -- 
    ack_4440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1966_delayed_1_0_1993_inst_ack_1, ack => convolve_CP_4061_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	112 
    -- CP-element group 121: 	120 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_sample_start_
      -- 
    rr_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(121), ack => type_cast_1999_inst_req_0); -- 
    convolve_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(112) & convolve_CP_4061_elements(120) & convolve_CP_4061_elements(123);
      gj_convolve_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: 	126 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_update_start_
      -- 
    cr_4453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(122), ack => type_cast_1999_inst_req_1); -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(124) & convolve_CP_4061_elements(126);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Sample/ra
      -- CP-element group 123: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_sample_completed_
      -- 
    ra_4449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_0, ack => convolve_CP_4061_elements(123)); -- 
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_1999_update_completed_
      -- 
    ca_4454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_1, ack => convolve_CP_4061_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: 	120 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	138 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Sample/req
      -- 
    req_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(125), ack => WPIPE_maxpool_output_pipe_1997_inst_req_0); -- 
    convolve_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(124) & convolve_CP_4061_elements(120) & convolve_CP_4061_elements(138) & convolve_CP_4061_elements(127);
      gj_convolve_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	122 
    -- CP-element group 126: 	118 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Update/req
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Sample/ack
      -- 
    ack_4463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1997_inst_ack_0, ack => convolve_CP_4061_elements(126)); -- 
    req_4467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(126), ack => WPIPE_maxpool_output_pipe_1997_inst_req_1); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	136 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_1997_Update/ack
      -- 
    ack_4468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1997_inst_ack_1, ack => convolve_CP_4061_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	30 
    -- CP-element group 128: 	95 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Sample/req
      -- CP-element group 128: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Sample/$entry
      -- 
    req_4476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(128), ack => W_next_sum_1971_delayed_1_0_2001_inst_req_0); -- 
    convolve_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(30) & convolve_CP_4061_elements(95) & convolve_CP_4061_elements(130);
      gj_convolve_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	134 
    -- CP-element group 129: 	137 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Update/req
      -- CP-element group 129: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_update_start_
      -- 
    req_4481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(129), ack => W_next_sum_1971_delayed_1_0_2001_inst_req_1); -- 
    convolve_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(134) & convolve_CP_4061_elements(137) & convolve_CP_4061_elements(131);
      gj_convolve_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	26 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	93 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Sample/ack
      -- CP-element group 130: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Sample/$exit
      -- 
    ack_4477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1971_delayed_1_0_2001_inst_ack_0, ack => convolve_CP_4061_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	136 
    -- CP-element group 131: 	132 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_Update/ack
      -- CP-element group 131: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/assign_stmt_2003_update_completed_
      -- 
    ack_4482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1971_delayed_1_0_2001_inst_ack_1, ack => convolve_CP_4061_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: 	116 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_sample_start_
      -- 
    rr_4490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(132), ack => type_cast_2007_inst_req_0); -- 
    convolve_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(131) & convolve_CP_4061_elements(116) & convolve_CP_4061_elements(134);
      gj_convolve_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	137 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Update/cr
      -- CP-element group 133: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_update_start_
      -- 
    cr_4495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(133), ack => type_cast_2007_inst_req_1); -- 
    convolve_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(135) & convolve_CP_4061_elements(137);
      gj_convolve_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	129 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	114 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Sample/$exit
      -- 
    ra_4491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2007_inst_ack_0, ack => convolve_CP_4061_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/type_cast_2007_Update/ca
      -- 
    ca_4496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2007_inst_ack_1, ack => convolve_CP_4061_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: 	127 
    -- CP-element group 136: 	131 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Sample/$entry
      -- 
    req_4504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(136), ack => WPIPE_maxpool_output_pipe_2005_inst_req_0); -- 
    convolve_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(135) & convolve_CP_4061_elements(127) & convolve_CP_4061_elements(131) & convolve_CP_4061_elements(138);
      gj_convolve_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	129 
    -- CP-element group 137: 	133 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Update/req
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Sample/$exit
      -- 
    ack_4505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2005_inst_ack_0, ack => convolve_CP_4061_elements(137)); -- 
    req_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(137), ack => WPIPE_maxpool_output_pipe_2005_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	125 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_Update/ack
      -- CP-element group 138: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/WPIPE_maxpool_output_pipe_2005_update_completed_
      -- 
    ack_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2005_inst_ack_1, ack => convolve_CP_4061_elements(138)); -- 
    -- CP-element group 139:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	19 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	20 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4061_elements(139) is a control-delay.
    cp_element_139_delay: control_delay_element  generic map(name => " 139_delay", delay_value => 1)  port map(req => convolve_CP_4061_elements(19), ack => convolve_CP_4061_elements(139), clk => clk, reset =>reset);
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	108 
    -- CP-element group 140: 	102 
    -- CP-element group 140: 	105 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	16 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_1833/do_while_stmt_1858/do_while_stmt_1858_loop_body/$exit
      -- 
    convolve_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4061_elements(138) & convolve_CP_4061_elements(108) & convolve_CP_4061_elements(102) & convolve_CP_4061_elements(105);
      gj_convolve_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4061_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	15 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_exit/$exit
      -- CP-element group 141: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_exit/ack
      -- 
    ack_4515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1858_branch_ack_0, ack => convolve_CP_4061_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	15 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_taken/$exit
      -- CP-element group 142: 	 branch_block_stmt_1833/do_while_stmt_1858/loop_taken/ack
      -- 
    ack_4519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1858_branch_ack_1, ack => convolve_CP_4061_elements(142)); -- 
    -- CP-element group 143:  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	13 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	2 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1833/do_while_stmt_1858/$exit
      -- 
    convolve_CP_4061_elements(143) <= convolve_CP_4061_elements(13);
    -- CP-element group 144:  merge  fork  transition  place  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	0 
    -- CP-element group 144: 	2 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	10 
    -- CP-element group 144: 	8 
    -- CP-element group 144: 	5 
    -- CP-element group 144: 	3 
    -- CP-element group 144:  members (19) 
      -- CP-element group 144: 	 branch_block_stmt_1833/merge_stmt_1834_PhiAck/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/merge_stmt_1834_PhiAck/$exit
      -- CP-element group 144: 	 branch_block_stmt_1833/merge_stmt_1834__exit__
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857__entry__
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1833/merge_stmt_1834_PhiAck/dummy
      -- CP-element group 144: 	 branch_block_stmt_1833/merge_stmt_1834_PhiReqMerge
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_num_out_pipe_1836_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/RPIPE_size_pipe_1839_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1843_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1833/assign_stmt_1837_to_assign_stmt_1857/slice_1847_Update/cr
      -- 
    rr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(144), ack => RPIPE_num_out_pipe_1836_inst_req_0); -- 
    rr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(144), ack => RPIPE_size_pipe_1839_inst_req_0); -- 
    cr_4119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(144), ack => slice_1843_inst_req_1); -- 
    cr_4133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4061_elements(144), ack => slice_1847_inst_req_1); -- 
    convolve_CP_4061_elements(144) <= OrReduce(convolve_CP_4061_elements(0) & convolve_CP_4061_elements(2));
    convolve_do_while_stmt_1858_terminator_4520: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1858_terminator_4520", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4061_elements(16),loop_continue => convolve_CP_4061_elements(142),loop_terminate => convolve_CP_4061_elements(141),loop_back => convolve_CP_4061_elements(14),loop_exit => convolve_CP_4061_elements(13),clk => clk, reset => reset); -- 
    phi_stmt_1860_phi_seq_4198_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4061_elements(33);
      convolve_CP_4061_elements(36)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4061_elements(36);
      convolve_CP_4061_elements(37)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4061_elements(38);
      convolve_CP_4061_elements(34) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4061_elements(31);
      convolve_CP_4061_elements(40)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4061_elements(42);
      convolve_CP_4061_elements(41)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4061_elements(43);
      convolve_CP_4061_elements(32) <= phi_mux_reqs(1);
      phi_stmt_1860_phi_seq_4198 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1860_phi_seq_4198") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4061_elements(27), 
          phi_sample_ack => convolve_CP_4061_elements(28), 
          phi_update_req => convolve_CP_4061_elements(29), 
          phi_update_ack => convolve_CP_4061_elements(30), 
          phi_mux_ack => convolve_CP_4061_elements(35), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1864_phi_seq_4242_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4061_elements(52);
      convolve_CP_4061_elements(55)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4061_elements(55);
      convolve_CP_4061_elements(56)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4061_elements(57);
      convolve_CP_4061_elements(53) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4061_elements(50);
      convolve_CP_4061_elements(59)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4061_elements(61);
      convolve_CP_4061_elements(60)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4061_elements(62);
      convolve_CP_4061_elements(51) <= phi_mux_reqs(1);
      phi_stmt_1864_phi_seq_4242 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1864_phi_seq_4242") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4061_elements(46), 
          phi_sample_ack => convolve_CP_4061_elements(47), 
          phi_update_req => convolve_CP_4061_elements(48), 
          phi_update_ack => convolve_CP_4061_elements(49), 
          phi_mux_ack => convolve_CP_4061_elements(54), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1868_phi_seq_4286_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4061_elements(67);
      convolve_CP_4061_elements(72)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4061_elements(74);
      convolve_CP_4061_elements(73)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4061_elements(75);
      convolve_CP_4061_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4061_elements(69);
      convolve_CP_4061_elements(76)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4061_elements(76);
      convolve_CP_4061_elements(77)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4061_elements(78);
      convolve_CP_4061_elements(70) <= phi_mux_reqs(1);
      phi_stmt_1868_phi_seq_4286 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1868_phi_seq_4286") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4061_elements(21), 
          phi_sample_ack => convolve_CP_4061_elements(65), 
          phi_update_req => convolve_CP_4061_elements(23), 
          phi_update_ack => convolve_CP_4061_elements(66), 
          phi_mux_ack => convolve_CP_4061_elements(71), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4150_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4061_elements(17);
        preds(1)  <= convolve_CP_4061_elements(18);
        entry_tmerge_4150 : transition_merge -- 
          generic map(name => " entry_tmerge_4150")
          port map (preds => preds, symbol_out => convolve_CP_4061_elements(19));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1971_wire : std_logic_vector(15 downto 0);
    signal ADD_u31_u31_1932_wire : std_logic_vector(30 downto 0);
    signal MUX_1972_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1920_1920_delayed_1_0_1943 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1946_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1952_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2011_wire : std_logic_vector(0 downto 0);
    signal SUB_u31_u31_1887_1887_delayed_1_0_1908 : std_logic_vector(30 downto 0);
    signal acc_1864 : std_logic_vector(15 downto 0);
    signal acc_val_1920 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1992 : std_logic_vector(7 downto 0);
    signal acc_val_up_1988 : std_logic_vector(7 downto 0);
    signal acc_var_1857 : std_logic_vector(15 downto 0);
    signal all_done_flag_1980 : std_logic_vector(0 downto 0);
    signal iread_1876 : std_logic_vector(15 downto 0);
    signal ival_1880 : std_logic_vector(15 downto 0);
    signal konst_1906_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1923_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1929_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1931_wire_constant : std_logic_vector(30 downto 0);
    signal konst_1970_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1983_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1894 : std_logic_vector(15 downto 0);
    signal kval_1898 : std_logic_vector(15 downto 0);
    signal mcount_var_1852 : std_logic_vector(30 downto 0);
    signal mul_val_1903 : std_logic_vector(15 downto 0);
    signal mycount_1860 : std_logic_vector(30 downto 0);
    signal n_out_count_1975 : std_logic_vector(15 downto 0);
    signal n_out_count_1975_1870_buffered : std_logic_vector(15 downto 0);
    signal nacc_1926 : std_logic_vector(15 downto 0);
    signal nacc_1926_1867_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1913 : std_logic_vector(0 downto 0);
    signal next_sum_1966_delayed_1_0_1995 : std_logic_vector(0 downto 0);
    signal next_sum_1971_delayed_1_0_2003 : std_logic_vector(0 downto 0);
    signal nmycount_1934 : std_logic_vector(30 downto 0);
    signal nmycount_1934_1863_buffered : std_logic_vector(30 downto 0);
    signal num_out_1837 : std_logic_vector(15 downto 0);
    signal out_count_1868 : std_logic_vector(15 downto 0);
    signal out_done_flag_1939 : std_logic_vector(0 downto 0);
    signal pingpong_1844 : std_logic_vector(0 downto 0);
    signal send_back1_1949 : std_logic_vector(0 downto 0);
    signal send_back2_1955 : std_logic_vector(0 downto 0);
    signal size_1848 : std_logic_vector(30 downto 0);
    signal size_read_1840 : std_logic_vector(31 downto 0);
    signal temp1_1884 : std_logic_vector(15 downto 0);
    signal temp2_1888 : std_logic_vector(15 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1916_wire : std_logic_vector(15 downto 0);
    signal type_cast_1918_wire : std_logic_vector(15 downto 0);
    signal type_cast_1968_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1999_wire : std_logic_vector(7 downto 0);
    signal type_cast_2007_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1857 <= "0000000000000000";
    konst_1906_wire_constant <= "0000000000000000000000000000001";
    konst_1923_wire_constant <= "0000000000000000";
    konst_1929_wire_constant <= "0000000000000000000000000000000";
    konst_1931_wire_constant <= "0000000000000000000000000000001";
    konst_1970_wire_constant <= "0000000000000001";
    konst_1983_wire_constant <= "1";
    mcount_var_1852 <= "0000000000000000000000000000000";
    type_cast_1872_wire_constant <= "0000000000000001";
    type_cast_1968_wire_constant <= "0000000000000001";
    phi_stmt_1860: Block -- phi operator 
      signal idata: std_logic_vector(61 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1852 & nmycount_1934_1863_buffered;
      req <= phi_stmt_1860_req_0 & phi_stmt_1860_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1860",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 31) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1860_ack_0,
          idata => idata,
          odata => mycount_1860,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1860
    phi_stmt_1864: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= acc_var_1857 & nacc_1926_1867_buffered;
      req <= phi_stmt_1864_req_0 & phi_stmt_1864_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1864",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1864_ack_0,
          idata => idata,
          odata => acc_1864,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1864
    phi_stmt_1868: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_out_count_1975_1870_buffered & type_cast_1872_wire_constant;
      req <= phi_stmt_1868_req_0 & phi_stmt_1868_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1868",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1868_ack_0,
          idata => idata,
          odata => out_count_1868,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1868
    -- flow-through select operator MUX_1893_inst
    kread_1894 <= temp2_1888 when (pingpong_1844(0) /=  '0') else temp1_1884;
    -- flow-through select operator MUX_1925_inst
    nacc_1926 <= konst_1923_wire_constant when (next_sum_1913(0) /=  '0') else acc_val_1920;
    -- flow-through select operator MUX_1933_inst
    nmycount_1934 <= konst_1929_wire_constant when (next_sum_1913(0) /=  '0') else ADD_u31_u31_1932_wire;
    -- flow-through select operator MUX_1972_inst
    MUX_1972_wire <= type_cast_1968_wire_constant when (out_done_flag_1939(0) /=  '0') else ADD_u16_u16_1971_wire;
    -- flow-through select operator MUX_1974_inst
    n_out_count_1975 <= MUX_1972_wire when (next_sum_1913(0) /=  '0') else out_count_1868;
    slice_1843_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1843_inst_req_0;
      slice_1843_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1843_inst_req_1;
      slice_1843_inst_ack_1<= update_ack(0);
      slice_1843_inst: SliceSplitProtocol generic map(name => "slice_1843_inst", in_data_width => 32, high_index => 31, low_index => 31, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => size_read_1840, dout => pingpong_1844, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1847_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1847_inst_req_0;
      slice_1847_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1847_inst_req_1;
      slice_1847_inst_ack_1<= update_ack(0);
      slice_1847_inst: SliceSplitProtocol generic map(name => "slice_1847_inst", in_data_width => 32, high_index => 30, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => size_read_1840, dout => size_1848, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1987_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1987_inst_req_0;
      slice_1987_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1987_inst_req_1;
      slice_1987_inst_ack_1<= update_ack(0);
      slice_1987_inst: SliceSplitProtocol generic map(name => "slice_1987_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1920, dout => acc_val_up_1988, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1991_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1991_inst_req_0;
      slice_1991_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1991_inst_req_1;
      slice_1991_inst_ack_1<= update_ack(0);
      slice_1991_inst: SliceSplitProtocol generic map(name => "slice_1991_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1920, dout => acc_val_dn_1992, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1966_delayed_1_0_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1966_delayed_1_0_1993_inst_req_0;
      W_next_sum_1966_delayed_1_0_1993_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1966_delayed_1_0_1993_inst_req_1;
      W_next_sum_1966_delayed_1_0_1993_inst_ack_1<= rack(0);
      W_next_sum_1966_delayed_1_0_1993_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1966_delayed_1_0_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1966_delayed_1_0_1995,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1971_delayed_1_0_2001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1971_delayed_1_0_2001_inst_req_0;
      W_next_sum_1971_delayed_1_0_2001_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1971_delayed_1_0_2001_inst_req_1;
      W_next_sum_1971_delayed_1_0_2001_inst_ack_1<= rack(0);
      W_next_sum_1971_delayed_1_0_2001_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1971_delayed_1_0_2001_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1971_delayed_1_0_2003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1975_1870_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1975_1870_buf_req_0;
      n_out_count_1975_1870_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1975_1870_buf_req_1;
      n_out_count_1975_1870_buf_ack_1<= rack(0);
      n_out_count_1975_1870_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1975_1870_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1975,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1975_1870_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1926_1867_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1926_1867_buf_req_0;
      nacc_1926_1867_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1926_1867_buf_req_1;
      nacc_1926_1867_buf_ack_1<= rack(0);
      nacc_1926_1867_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1926_1867_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1926_1867_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1934_1863_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1934_1863_buf_req_0;
      nmycount_1934_1863_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1934_1863_buf_req_1;
      nmycount_1934_1863_buf_ack_1<= rack(0);
      nmycount_1934_1863_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1934_1863_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 31,
        out_data_width => 31,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1934,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1934_1863_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1879_inst
    process(iread_1876) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1876(15 downto 0);
      ival_1880 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1897_inst
    process(kread_1894) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1894(15 downto 0);
      kval_1898 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1916_inst
    process(acc_1864) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1864(15 downto 0);
      type_cast_1916_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1918_inst
    process(mul_val_1903) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1903(15 downto 0);
      type_cast_1918_wire <= tmp_var; -- 
    end process;
    type_cast_1999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1999_inst_req_0;
      type_cast_1999_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1999_inst_req_1;
      type_cast_1999_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1966_delayed_1_0_1995(0);
      type_cast_1999_inst_gI: SplitGuardInterface generic map(name => "type_cast_1999_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1988,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_2007_inst_req_0;
      type_cast_2007_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_2007_inst_req_1;
      type_cast_2007_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1971_delayed_1_0_2003(0);
      type_cast_2007_inst_gI: SplitGuardInterface generic map(name => "type_cast_2007_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_2007_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1992,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2007_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1858_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2011_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1858_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1858_branch_req_0,
          ack0 => do_while_stmt_1858_branch_ack_0,
          ack1 => do_while_stmt_1858_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1919_inst
    process(type_cast_1916_wire, type_cast_1918_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1916_wire, type_cast_1918_wire, tmp_var);
      acc_val_1920 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1971_inst
    process(out_count_1868) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1868, konst_1970_wire_constant, tmp_var);
      ADD_u16_u16_1971_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u31_u31_1932_inst
    process(mycount_1860) -- 
      variable tmp_var : std_logic_vector(30 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1860, konst_1931_wire_constant, tmp_var);
      ADD_u31_u31_1932_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1948_inst
    process(NOT_u1_u1_1946_wire, NOT_u1_u1_1920_1920_delayed_1_0_1943) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1946_wire, NOT_u1_u1_1920_1920_delayed_1_0_1943, tmp_var);
      send_back1_1949 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1954_inst
    process(NOT_u1_u1_1952_wire, pingpong_1844) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1952_wire, pingpong_1844, tmp_var);
      send_back2_1955 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1979_inst
    process(out_done_flag_1939, next_sum_1913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1939, next_sum_1913, tmp_var);
      all_done_flag_1980 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1938_inst
    process(out_count_1868, num_out_1837) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1868, num_out_1837, tmp_var);
      out_done_flag_1939 <= tmp_var; --
    end process;
    -- binary operator EQ_u31_u1_1912_inst
    process(mycount_1860, SUB_u31_u31_1887_1887_delayed_1_0_1908) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1860, SUB_u31_u31_1887_1887_delayed_1_0_1908, tmp_var);
      next_sum_1913 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1902_inst
    process(kval_1898, ival_1880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1898, ival_1880, tmp_var);
      mul_val_1903 <= tmp_var; --
    end process;
    -- shared split operator group (9) : NOT_u1_u1_1942_inst 
    ApIntNot_group_9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pingpong_1844;
      NOT_u1_u1_1920_1920_delayed_1_0_1943 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1942_inst_req_0;
      NOT_u1_u1_1942_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1942_inst_req_1;
      NOT_u1_u1_1942_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_9_gI: SplitGuardInterface generic map(name => "ApIntNot_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- unary operator NOT_u1_u1_1946_inst
    process(out_done_flag_1939) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", out_done_flag_1939, tmp_var);
      NOT_u1_u1_1946_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1952_inst
    process(out_done_flag_1939) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", out_done_flag_1939, tmp_var);
      NOT_u1_u1_1952_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2011_inst
    process(all_done_flag_1980) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_1980, tmp_var);
      NOT_u1_u1_2011_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (13) : SUB_u31_u31_1907_inst 
    ApIntSub_group_13: Block -- 
      signal data_in: std_logic_vector(30 downto 0);
      signal data_out: std_logic_vector(30 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1848;
      SUB_u31_u31_1887_1887_delayed_1_0_1908 <= data_out(30 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u31_u31_1907_inst_req_0;
      SUB_u31_u31_1907_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u31_u31_1907_inst_req_1;
      SUB_u31_u31_1907_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_13_gI: SplitGuardInterface generic map(name => "ApIntSub_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 31,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 31,
          constant_operand => "0000000000000000000000000000001",
          constant_width => 31,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared inport operator group (0) : RPIPE_input_pipe1_1875_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1875_inst_req_0;
      RPIPE_input_pipe1_1875_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1875_inst_req_1;
      RPIPE_input_pipe1_1875_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1876 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1883_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1883_inst_req_0;
      RPIPE_kernel_pipe1_1883_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1883_inst_req_1;
      RPIPE_kernel_pipe1_1883_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not pingpong_1844(0);
      temp1_1884 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_kernel_pipe2_1887_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_1887_inst_req_0;
      RPIPE_kernel_pipe2_1887_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_1887_inst_req_1;
      RPIPE_kernel_pipe2_1887_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pingpong_1844(0);
      temp2_1888 <= data_out(15 downto 0);
      kernel_pipe2_read_2_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_2: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_num_out_pipe_1836_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1836_inst_req_0;
      RPIPE_num_out_pipe_1836_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1836_inst_req_1;
      RPIPE_num_out_pipe_1836_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1837 <= data_out(15 downto 0);
      num_out_pipe_read_3_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_3: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_size_pipe_1839_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1839_inst_req_0;
      RPIPE_size_pipe_1839_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1839_inst_req_1;
      RPIPE_size_pipe_1839_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_read_1840 <= data_out(31 downto 0);
      size_pipe_read_4_gI: SplitGuardInterface generic map(name => "size_pipe_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_4: InputPortRevised -- 
        generic map ( name => "size_pipe_read_4", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1982_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1982_inst_req_0;
      WPIPE_input_done_pipe_1982_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1982_inst_req_1;
      WPIPE_input_done_pipe_1982_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1980(0);
      data_in <= konst_1983_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1957_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1957_inst_req_0;
      WPIPE_kernel_pipe1_1957_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1957_inst_req_1;
      WPIPE_kernel_pipe1_1957_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_back1_1949(0);
      data_in <= kread_1894;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe2_1961_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_1961_inst_req_0;
      WPIPE_kernel_pipe2_1961_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_1961_inst_req_1;
      WPIPE_kernel_pipe2_1961_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_back2_1955(0);
      data_in <= kread_1894;
      kernel_pipe2_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_maxpool_output_pipe_1997_inst WPIPE_maxpool_output_pipe_2005_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1997_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2005_inst_req_0;
      WPIPE_maxpool_output_pipe_1997_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2005_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1997_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2005_inst_req_1;
      WPIPE_maxpool_output_pipe_1997_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2005_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1971_delayed_1_0_2003(0);
      guard_vector(1)  <= next_sum_1966_delayed_1_0_1995(0);
      data_in <= type_cast_1999_wire & type_cast_2007_wire;
      maxpool_output_pipe_write_3_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    pp : in  std_logic_vector(7 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 136)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  signal pp_buffer :  std_logic_vector(7 downto 0);
  signal pp_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_671_start: Boolean;
  signal loadKernelChannel_CP_671_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_fn_403_delayed_7_0_415_inst_req_1 : boolean;
  signal nfetch_val_434_369_buf_req_0 : boolean;
  signal CONCAT_u1_u32_449_inst_req_1 : boolean;
  signal WPIPE_size_pipe_442_inst_ack_0 : boolean;
  signal W_fn_403_delayed_7_0_415_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_392_inst_req_0 : boolean;
  signal nfetch_val_434_369_buf_req_1 : boolean;
  signal W_fetch_val_411_delayed_13_0_426_inst_req_1 : boolean;
  signal ptr_deref_421_load_0_ack_0 : boolean;
  signal CONCAT_u1_u32_449_inst_ack_1 : boolean;
  signal my_fetch_349_368_buf_ack_1 : boolean;
  signal W_fetch_val_411_delayed_13_0_426_inst_ack_1 : boolean;
  signal nfetch_val_434_369_buf_ack_1 : boolean;
  signal array_obj_ref_412_index_offset_req_1 : boolean;
  signal array_obj_ref_412_index_offset_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_396_inst_ack_1 : boolean;
  signal array_obj_ref_412_index_offset_req_0 : boolean;
  signal WPIPE_size_pipe_442_inst_req_1 : boolean;
  signal ptr_deref_421_load_0_req_1 : boolean;
  signal array_obj_ref_412_index_offset_ack_0 : boolean;
  signal WPIPE_size_pipe_442_inst_ack_1 : boolean;
  signal phi_stmt_366_req_0 : boolean;
  signal do_while_stmt_360_branch_ack_0 : boolean;
  signal W_fn_403_delayed_7_0_415_inst_req_0 : boolean;
  signal ptr_deref_421_load_0_ack_1 : boolean;
  signal phi_stmt_366_req_1 : boolean;
  signal W_fetch_val_411_delayed_13_0_426_inst_ack_0 : boolean;
  signal W_fn_403_delayed_7_0_415_inst_ack_0 : boolean;
  signal my_fetch_349_368_buf_req_1 : boolean;
  signal W_fn_409_delayed_13_0_423_inst_req_0 : boolean;
  signal nfetch_val_434_369_buf_ack_0 : boolean;
  signal W_fn_409_delayed_13_0_423_inst_ack_0 : boolean;
  signal addr_of_413_final_reg_req_0 : boolean;
  signal WPIPE_kernel_pipe2_396_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_392_inst_ack_0 : boolean;
  signal addr_of_413_final_reg_ack_0 : boolean;
  signal W_fn_409_delayed_13_0_423_inst_req_1 : boolean;
  signal W_fn_409_delayed_13_0_423_inst_ack_1 : boolean;
  signal phi_stmt_366_ack_0 : boolean;
  signal W_fetch_val_411_delayed_13_0_426_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_396_inst_ack_0 : boolean;
  signal addr_of_413_final_reg_req_1 : boolean;
  signal ptr_deref_421_load_0_req_0 : boolean;
  signal addr_of_413_final_reg_ack_1 : boolean;
  signal CONCAT_u1_u32_449_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_396_inst_req_0 : boolean;
  signal WPIPE_size_pipe_442_inst_req_0 : boolean;
  signal CONCAT_u1_u32_449_inst_ack_0 : boolean;
  signal my_fetch_349_368_buf_req_0 : boolean;
  signal my_fetch_349_368_buf_ack_0 : boolean;
  signal start_add_365_buf_ack_1 : boolean;
  signal array_obj_ref_343_index_offset_req_0 : boolean;
  signal array_obj_ref_343_index_offset_ack_0 : boolean;
  signal array_obj_ref_343_index_offset_req_1 : boolean;
  signal array_obj_ref_343_index_offset_ack_1 : boolean;
  signal do_while_stmt_360_branch_ack_1 : boolean;
  signal addr_of_344_final_reg_req_0 : boolean;
  signal addr_of_344_final_reg_ack_0 : boolean;
  signal addr_of_344_final_reg_req_1 : boolean;
  signal addr_of_344_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_392_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_392_inst_req_1 : boolean;
  signal start_add_365_buf_req_1 : boolean;
  signal ptr_deref_348_load_0_req_0 : boolean;
  signal ptr_deref_348_load_0_ack_0 : boolean;
  signal ptr_deref_348_load_0_req_1 : boolean;
  signal ptr_deref_348_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_357_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_357_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_357_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_357_inst_ack_1 : boolean;
  signal do_while_stmt_360_branch_req_0 : boolean;
  signal phi_stmt_362_req_0 : boolean;
  signal phi_stmt_362_req_1 : boolean;
  signal phi_stmt_362_ack_0 : boolean;
  signal nmycount_384_364_buf_req_0 : boolean;
  signal nmycount_384_364_buf_ack_0 : boolean;
  signal nmycount_384_364_buf_req_1 : boolean;
  signal nmycount_384_364_buf_ack_1 : boolean;
  signal start_add_365_buf_req_0 : boolean;
  signal start_add_365_buf_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 136) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(135 downto 128) <= pp;
  pp_buffer <= in_buffer_data_out(135 downto 128);
  in_buffer_data_in(tag_length + 135 downto 136) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 135 downto 136);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_671_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_671: Block -- control-path 
    signal loadKernelChannel_CP_671_elements: BooleanArray(97 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_671_elements(0) <= loadKernelChannel_CP_671_start;
    loadKernelChannel_CP_671_symbol <= loadKernelChannel_CP_671_elements(97);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_update_start_
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_resized_1
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_computed_1
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_complete/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_complete/req
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_update_start_
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_sample_start_
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Sample/rr
      -- 
    rr_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => RPIPE_input_done_pipe_357_inst_req_0); -- 
    req_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_343_index_offset_req_0); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_343_index_offset_req_1); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => addr_of_344_final_reg_req_1); -- 
    cr_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => ptr_deref_348_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Sample/ack
      -- 
    ack_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_343_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_sample_start_
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_offset_calculated
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/array_obj_ref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_request/$entry
      -- CP-element group 2: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_request/req
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_343_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(2)); -- 
    req_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(2), ack => addr_of_344_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_sample_completed_
      -- CP-element group 3: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_request/$exit
      -- CP-element group 3: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_request/ack
      -- 
    ack_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_344_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_update_completed_
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_complete/$exit
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/addr_of_344_complete/ack
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_sample_start_
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_address_resized
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/word_0/rr
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_344_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(4)); -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(4), ack => ptr_deref_348_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_sample_completed_
      -- CP-element group 5: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Sample/word_access_start/word_0/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_348_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_update_completed_
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/$exit
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/ptr_deref_348_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/ptr_deref_348_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/ptr_deref_348_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_334_to_assign_stmt_358/ptr_deref_348_Update/ptr_deref_348_Merge/merge_ack
      -- 
    ca_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_348_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_sample_completed_
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_update_start_
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Sample/ra
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Update/$entry
      -- CP-element group 7: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Update/cr
      -- 
    ra_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_357_inst_ack_0, ack => loadKernelChannel_CP_671_elements(7)); -- 
    cr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(7), ack => RPIPE_input_done_pipe_357_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_update_completed_
      -- CP-element group 8: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Update/$exit
      -- CP-element group 8: 	 assign_stmt_334_to_assign_stmt_358/RPIPE_input_done_pipe_357_Update/ca
      -- 
    ca_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_357_inst_ack_1, ack => loadKernelChannel_CP_671_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_334_to_assign_stmt_358/$exit
      -- CP-element group 9: 	 branch_block_stmt_359/$entry
      -- CP-element group 9: 	 branch_block_stmt_359/branch_block_stmt_359__entry__
      -- CP-element group 9: 	 branch_block_stmt_359/do_while_stmt_360__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(6) & loadKernelChannel_CP_671_elements(8) & loadKernelChannel_CP_671_elements(1);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	93 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	94 
    -- CP-element group 10: 	95 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_Update/cr
      -- CP-element group 10: 	 assign_stmt_450/$entry
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_Update/$entry
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_update_start_
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_359/$exit
      -- CP-element group 10: 	 branch_block_stmt_359/branch_block_stmt_359__exit__
      -- CP-element group 10: 	 branch_block_stmt_359/do_while_stmt_360__exit__
      -- CP-element group 10: 	 assign_stmt_450/CONCAT_u1_u32_449_sample_start_
      -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => CONCAT_u1_u32_449_inst_req_1); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => CONCAT_u1_u32_449_inst_req_0); -- 
    loadKernelChannel_CP_671_elements(10) <= loadKernelChannel_CP_671_elements(93);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_359/do_while_stmt_360/$entry
      -- CP-element group 11: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360__entry__
      -- 
    loadKernelChannel_CP_671_elements(11) <= loadKernelChannel_CP_671_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	93 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360__exit__
      -- 
    -- Element group loadKernelChannel_CP_671_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_359/do_while_stmt_360/loop_back
      -- 
    -- Element group loadKernelChannel_CP_671_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	91 
    -- CP-element group 14: 	92 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_359/do_while_stmt_360/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_359/do_while_stmt_360/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_359/do_while_stmt_360/condition_done
      -- 
    loadKernelChannel_CP_671_elements(14) <= loadKernelChannel_CP_671_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	90 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_359/do_while_stmt_360/loop_body_done
      -- 
    loadKernelChannel_CP_671_elements(15) <= loadKernelChannel_CP_671_elements(90);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_671_elements(16) <= loadKernelChannel_CP_671_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	30 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_671_elements(17) <= loadKernelChannel_CP_671_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	68 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	67 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	89 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	89 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/condition_evaluated
      -- 
    condition_evaluated_808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(19), ack => do_while_stmt_360_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(23) & loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(89);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(24) & loadKernelChannel_CP_671_elements(41) & loadKernelChannel_CP_671_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	82 
    -- CP-element group 21: 	78 
    -- CP-element group 21: 	86 
    -- CP-element group 21: 	90 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(26) & loadKernelChannel_CP_671_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(25) & loadKernelChannel_CP_671_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	69 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	83 
    -- CP-element group 25: 	75 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(69) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(64) & loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(83) & loadKernelChannel_CP_671_elements(75);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	69 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	81 
    -- CP-element group 27: 	73 
    -- CP-element group 27: 	60 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_update_completed__ps
      -- 
    req_974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(27), ack => array_obj_ref_412_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(28) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_loopback_sample_req_ps
      -- 
    phi_stmt_362_loopback_sample_req_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_362_loopback_sample_req_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(29), ack => phi_stmt_362_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(30) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_entry_sample_req_ps
      -- 
    phi_stmt_362_entry_sample_req_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_362_entry_sample_req_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(31), ack => phi_stmt_362_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_362_phi_mux_ack_ps
      -- 
    phi_stmt_362_phi_mux_ack_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_362_ack_0, ack => loadKernelChannel_CP_671_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Sample/req
      -- 
    req_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(33), ack => nmycount_384_364_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_update_start_
      -- CP-element group 34: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Update/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(34), ack => nmycount_384_364_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Sample/ack
      -- 
    ack_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_384_364_buf_ack_0, ack => loadKernelChannel_CP_671_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nmycount_364_Update/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_384_364_buf_ack_1, ack => loadKernelChannel_CP_671_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Sample/req
      -- 
    req_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(37), ack => start_add_365_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Update/req
      -- CP-element group 38: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_update_start_
      -- CP-element group 38: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Update/$entry
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(38), ack => start_add_365_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Sample/ack
      -- 
    ack_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_365_buf_ack_0, ack => loadKernelChannel_CP_671_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_start_add_365_update_completed_
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_365_buf_ack_1, ack => loadKernelChannel_CP_671_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	80 
    -- CP-element group 41: 	84 
    -- CP-element group 41: 	88 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(80) & loadKernelChannel_CP_671_elements(84) & loadKernelChannel_CP_671_elements(88);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	87 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(64) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(87);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_sample_start__ps
      -- 
    loadKernelChannel_CP_671_elements(43) <= loadKernelChannel_CP_671_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_update_start__ps
      -- 
    loadKernelChannel_CP_671_elements(45) <= loadKernelChannel_CP_671_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	85 
    -- CP-element group 46: 	60 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_671_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(47) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_loopback_sample_req
      -- 
    phi_stmt_366_loopback_sample_req_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_366_loopback_sample_req_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(48), ack => phi_stmt_366_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(49) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_entry_sample_req_ps
      -- 
    phi_stmt_366_entry_sample_req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_366_entry_sample_req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(50), ack => phi_stmt_366_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/phi_stmt_366_phi_mux_ack_ps
      -- 
    phi_stmt_366_phi_mux_ack_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_366_ack_0, ack => loadKernelChannel_CP_671_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Sample/req
      -- 
    req_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(52), ack => my_fetch_349_368_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Update/req
      -- CP-element group 53: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_update_start_
      -- CP-element group 53: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Update/$entry
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(53), ack => my_fetch_349_368_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Sample/ack
      -- 
    ack_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_349_368_buf_ack_0, ack => loadKernelChannel_CP_671_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_my_fetch_368_Update/$exit
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_349_368_buf_ack_1, ack => loadKernelChannel_CP_671_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Sample/$entry
      -- 
    req_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(56), ack => nfetch_val_434_369_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Update/req
      -- CP-element group 57: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_update_start_
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(57), ack => nfetch_val_434_369_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Sample/$exit
      -- 
    ack_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_434_369_buf_ack_0, ack => loadKernelChannel_CP_671_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/R_nfetch_val_369_update_completed_
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_434_369_buf_ack_1, ack => loadKernelChannel_CP_671_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Sample/$entry
      -- 
    req_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(60), ack => WPIPE_kernel_pipe1_392_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_update_start_
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Update/req
      -- CP-element group 61: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Update/$entry
      -- 
    ack_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_392_inst_ack_0, ack => loadKernelChannel_CP_671_elements(61)); -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(61), ack => WPIPE_kernel_pipe1_392_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	90 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe1_392_Update/$exit
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_392_inst_ack_1, ack => loadKernelChannel_CP_671_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_sample_start_
      -- 
    req_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(63), ack => WPIPE_kernel_pipe2_396_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Update/req
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_update_start_
      -- CP-element group 64: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_sample_completed_
      -- 
    ack_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_396_inst_ack_0, ack => loadKernelChannel_CP_671_elements(64)); -- 
    req_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(64), ack => WPIPE_kernel_pipe2_396_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	90 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/WPIPE_kernel_pipe2_396_update_completed_
      -- 
    ack_949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_396_inst_ack_1, ack => loadKernelChannel_CP_671_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	70 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	71 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	71 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_request/$entry
      -- CP-element group 66: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_request/req
      -- 
    req_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(66), ack => addr_of_413_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(70) & loadKernelChannel_CP_671_elements(71);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	18 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	72 
    -- CP-element group 67: 	79 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	72 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_update_start_
      -- CP-element group 67: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_complete/$entry
      -- CP-element group 67: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_complete/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(67), ack => addr_of_413_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(72) & loadKernelChannel_CP_671_elements(79);
      gj_loadKernelChannel_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	18 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: 	71 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_update_start
      -- CP-element group 68: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Update/req
      -- CP-element group 68: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Update/$entry
      -- 
    req_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(68), ack => array_obj_ref_412_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(70) & loadKernelChannel_CP_671_elements(71);
      gj_loadKernelChannel_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	27 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	90 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	25 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_sample_complete
      -- 
    ack_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_412_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(69)); -- 
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (8) 
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_root_address_calculated
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_offset_calculated
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_final_index_sum_regn_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_base_plus_offset/$entry
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_base_plus_offset/$exit
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_base_plus_offset/sum_rename_req
      -- CP-element group 70: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/array_obj_ref_412_base_plus_offset/sum_rename_ack
      -- 
    ack_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_412_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	66 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	68 
    -- CP-element group 71: 	66 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_request/$exit
      -- CP-element group 71: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_request/ack
      -- 
    ack_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_413_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(71)); -- 
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	67 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	77 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	67 
    -- CP-element group 72:  members (19) 
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_plus_offset/$entry
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_plus_offset/sum_rename_req
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_plus_offset/sum_rename_ack
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_word_addrgen/root_register_req
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_word_addrgen/$entry
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_word_addrgen/$exit
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_word_addrgen/root_register_ack
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_addr_resize/base_resize_req
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_plus_offset/$exit
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_addr_resize/base_resize_ack
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/addr_of_413_complete/ack
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_addr_resize/$exit
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_addr_resize/$entry
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_address_resized
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_root_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_word_address_calculated
      -- CP-element group 72: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_base_address_calculated
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_413_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	27 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Sample/req
      -- CP-element group 73: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Sample/$entry
      -- 
    req_1003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(73), ack => W_fn_403_delayed_7_0_415_inst_req_0); -- 
    loadKernelChannel_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(75);
      gj_loadKernelChannel_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	79 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Update/req
      -- CP-element group 74: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_update_start_
      -- 
    req_1008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(74), ack => W_fn_403_delayed_7_0_415_inst_req_1); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(79) & loadKernelChannel_CP_671_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	25 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Sample/ack
      -- CP-element group 75: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Sample/$exit
      -- 
    ack_1004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_403_delayed_7_0_415_inst_ack_0, ack => loadKernelChannel_CP_671_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Update/ack
      -- CP-element group 76: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_417_update_completed_
      -- 
    ack_1009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_403_delayed_7_0_415_inst_ack_1, ack => loadKernelChannel_CP_671_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	72 
    -- CP-element group 77: 	76 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/word_0/$entry
      -- 
    rr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(77), ack => ptr_deref_421_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(72) & loadKernelChannel_CP_671_elements(76) & loadKernelChannel_CP_671_elements(79);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	21 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/$entry
      -- CP-element group 78: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/word_0/cr
      -- CP-element group 78: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_update_start_
      -- 
    cr_1053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(78), ack => ptr_deref_421_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	67 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/word_0/ra
      -- CP-element group 79: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Sample/word_access_start/word_0/$exit
      -- 
    ra_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_421_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(79)); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	90 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	41 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/ptr_deref_421_Merge/$entry
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/ptr_deref_421_Merge/$exit
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/ptr_deref_421_Merge/merge_req
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/ptr_deref_421_Update/ptr_deref_421_Merge/merge_ack
      -- 
    ca_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_421_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	27 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Sample/req
      -- CP-element group 81: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_sample_start_
      -- 
    req_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(81), ack => W_fn_409_delayed_13_0_423_inst_req_0); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	21 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_update_start_
      -- CP-element group 82: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Update/req
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(82), ack => W_fn_409_delayed_13_0_423_inst_req_1); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	25 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Sample/ack
      -- 
    ack_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_409_delayed_13_0_423_inst_ack_0, ack => loadKernelChannel_CP_671_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	90 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	41 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_425_Update/ack
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_409_delayed_13_0_423_inst_ack_1, ack => loadKernelChannel_CP_671_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	46 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Sample/req
      -- 
    req_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(85), ack => W_fetch_val_411_delayed_13_0_426_inst_req_0); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	21 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	88 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_update_start_
      -- CP-element group 86: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Update/req
      -- 
    req_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(86), ack => W_fetch_val_411_delayed_13_0_426_inst_req_1); -- 
    loadKernelChannel_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(88);
      gj_loadKernelChannel_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	42 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_sample_completed_
      -- 
    ack_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_411_delayed_13_0_426_inst_ack_0, ack => loadKernelChannel_CP_671_elements(87)); -- 
    -- CP-element group 88:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	41 
    -- CP-element group 88: 	86 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/assign_stmt_428_Update/ack
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_411_delayed_13_0_426_inst_ack_1, ack => loadKernelChannel_CP_671_elements(88)); -- 
    -- CP-element group 89:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	18 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	19 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_671_elements(18), ack => loadKernelChannel_CP_671_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  join  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	69 
    -- CP-element group 90: 	62 
    -- CP-element group 90: 	21 
    -- CP-element group 90: 	80 
    -- CP-element group 90: 	65 
    -- CP-element group 90: 	84 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	15 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_359/do_while_stmt_360/do_while_stmt_360_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(69) & loadKernelChannel_CP_671_elements(62) & loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(80) & loadKernelChannel_CP_671_elements(65) & loadKernelChannel_CP_671_elements(84) & loadKernelChannel_CP_671_elements(88);
      gj_loadKernelChannel_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	14 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_359/do_while_stmt_360/loop_exit/ack
      -- CP-element group 91: 	 branch_block_stmt_359/do_while_stmt_360/loop_exit/$exit
      -- 
    ack_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_360_branch_ack_0, ack => loadKernelChannel_CP_671_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	14 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_359/do_while_stmt_360/loop_taken/$exit
      -- CP-element group 92: 	 branch_block_stmt_359/do_while_stmt_360/loop_taken/ack
      -- 
    ack_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_360_branch_ack_1, ack => loadKernelChannel_CP_671_elements(92)); -- 
    -- CP-element group 93:  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	10 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_359/do_while_stmt_360/$exit
      -- 
    loadKernelChannel_CP_671_elements(93) <= loadKernelChannel_CP_671_elements(12);
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	10 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_450/CONCAT_u1_u32_449_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_450/CONCAT_u1_u32_449_Sample/ra
      -- CP-element group 94: 	 assign_stmt_450/CONCAT_u1_u32_449_sample_completed_
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_449_inst_ack_0, ack => loadKernelChannel_CP_671_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	10 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 assign_stmt_450/CONCAT_u1_u32_449_Update/ca
      -- CP-element group 95: 	 assign_stmt_450/CONCAT_u1_u32_449_Update/$exit
      -- CP-element group 95: 	 assign_stmt_450/WPIPE_size_pipe_442_sample_start_
      -- CP-element group 95: 	 assign_stmt_450/CONCAT_u1_u32_449_update_completed_
      -- CP-element group 95: 	 assign_stmt_450/WPIPE_size_pipe_442_Sample/$entry
      -- CP-element group 95: 	 assign_stmt_450/WPIPE_size_pipe_442_Sample/req
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u32_449_inst_ack_1, ack => loadKernelChannel_CP_671_elements(95)); -- 
    req_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(95), ack => WPIPE_size_pipe_442_inst_req_0); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_Sample/ack
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_Update/$entry
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_Update/req
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_Sample/$exit
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_sample_completed_
      -- CP-element group 96: 	 assign_stmt_450/WPIPE_size_pipe_442_update_start_
      -- 
    ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_442_inst_ack_0, ack => loadKernelChannel_CP_671_elements(96)); -- 
    req_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(96), ack => WPIPE_size_pipe_442_inst_req_1); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 assign_stmt_450/WPIPE_size_pipe_442_Update/$exit
      -- CP-element group 97: 	 assign_stmt_450/WPIPE_size_pipe_442_Update/ack
      -- CP-element group 97: 	 assign_stmt_450/$exit
      -- CP-element group 97: 	 assign_stmt_450/WPIPE_size_pipe_442_update_completed_
      -- CP-element group 97: 	 $exit
      -- 
    ack_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_442_inst_ack_1, ack => loadKernelChannel_CP_671_elements(97)); -- 
    loadKernelChannel_do_while_stmt_360_terminator_1097: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_360_terminator_1097", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_671_elements(15),loop_continue => loadKernelChannel_CP_671_elements(92),loop_terminate => loadKernelChannel_CP_671_elements(91),loop_back => loadKernelChannel_CP_671_elements(13),loop_exit => loadKernelChannel_CP_671_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_362_phi_seq_867_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(28);
      loadKernelChannel_CP_671_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(35);
      loadKernelChannel_CP_671_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(36);
      loadKernelChannel_CP_671_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(30);
      loadKernelChannel_CP_671_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(39);
      loadKernelChannel_CP_671_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(40);
      loadKernelChannel_CP_671_elements(31) <= phi_mux_reqs(1);
      phi_stmt_362_phi_seq_867 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_362_phi_seq_867") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(26), 
          phi_update_req => loadKernelChannel_CP_671_elements(22), 
          phi_update_ack => loadKernelChannel_CP_671_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_366_phi_seq_921_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(49);
      loadKernelChannel_CP_671_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(54);
      loadKernelChannel_CP_671_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(55);
      loadKernelChannel_CP_671_elements(50) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(47);
      loadKernelChannel_CP_671_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(58);
      loadKernelChannel_CP_671_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(59);
      loadKernelChannel_CP_671_elements(48) <= phi_mux_reqs(1);
      phi_stmt_366_phi_seq_921 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_366_phi_seq_921") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(44), 
          phi_update_req => loadKernelChannel_CP_671_elements(45), 
          phi_update_ack => loadKernelChannel_CP_671_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_809_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_671_elements(16);
        preds(1)  <= loadKernelChannel_CP_671_elements(17);
        entry_tmerge_809 : transition_merge -- 
          generic map(name => " entry_tmerge_809")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_671_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_375_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_402_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u1_u32_449_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_388_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_411_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_411_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_411_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_342_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_342_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_376_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_439_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_447_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_440_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_343_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_343_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_343_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_343_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_343_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_343_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_412_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_345 : std_logic_vector(31 downto 0);
    signal fetch_addr_414 : std_logic_vector(31 downto 0);
    signal fetch_val_366 : std_logic_vector(63 downto 0);
    signal fetch_val_411_delayed_13_0_428 : std_logic_vector(63 downto 0);
    signal first_fill_354 : std_logic_vector(0 downto 0);
    signal fn_403_delayed_7_0_417 : std_logic_vector(0 downto 0);
    signal fn_405 : std_logic_vector(0 downto 0);
    signal fn_409_delayed_13_0_425 : std_logic_vector(0 downto 0);
    signal fv_422 : std_logic_vector(63 downto 0);
    signal konst_332_wire_constant : std_logic_vector(63 downto 0);
    signal konst_352_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_374_wire_constant : std_logic_vector(63 downto 0);
    signal konst_377_wire_constant : std_logic_vector(63 downto 0);
    signal konst_382_wire_constant : std_logic_vector(63 downto 0);
    signal konst_401_wire_constant : std_logic_vector(63 downto 0);
    signal konst_403_wire_constant : std_logic_vector(63 downto 0);
    signal konst_410_wire_constant : std_logic_vector(63 downto 0);
    signal konst_438_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_349 : std_logic_vector(63 downto 0);
    signal my_fetch_349_368_buffered : std_logic_vector(63 downto 0);
    signal my_num1_379 : std_logic_vector(63 downto 0);
    signal mycount_362 : std_logic_vector(63 downto 0);
    signal nfetch_val_434 : std_logic_vector(63 downto 0);
    signal nfetch_val_434_369_buffered : std_logic_vector(63 downto 0);
    signal nmycount_384 : std_logic_vector(63 downto 0);
    signal nmycount_384_364_buffered : std_logic_vector(63 downto 0);
    signal pingpong_338 : std_logic_vector(0 downto 0);
    signal ptr_deref_348_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_348_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_348_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_348_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_348_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_421_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_421_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_421_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_421_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_421_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_334 : std_logic_vector(63 downto 0);
    signal start_add_365_buffered : std_logic_vector(63 downto 0);
    signal start_next_358 : std_logic_vector(0 downto 0);
    signal type_cast_448_wire : std_logic_vector(30 downto 0);
    signal var_val_390 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_343_constant_part_of_offset <= "00000000000000";
    array_obj_ref_343_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_343_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_343_resized_base_address <= "00000000000000";
    array_obj_ref_412_constant_part_of_offset <= "00000000000000";
    array_obj_ref_412_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_412_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_412_resized_base_address <= "00000000000000";
    konst_332_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_374_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_377_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_382_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_403_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_410_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_348_word_offset_0 <= "00000000000000";
    ptr_deref_421_word_offset_0 <= "00000000000000";
    phi_stmt_362: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_384_364_buffered & start_add_365_buffered;
      req <= phi_stmt_362_req_0 & phi_stmt_362_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_362",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_362_ack_0,
          idata => idata,
          odata => mycount_362,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_362
    phi_stmt_366: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch_349_368_buffered & nfetch_val_434_369_buffered;
      req <= phi_stmt_366_req_0 & phi_stmt_366_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_366",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_366_ack_0,
          idata => idata,
          odata => fetch_val_366,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_366
    -- flow-through select operator MUX_433_inst
    nfetch_val_434 <= fv_422 when (fn_409_delayed_13_0_425(0) /=  '0') else fetch_val_411_delayed_13_0_428;
    W_fetch_val_411_delayed_13_0_426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_411_delayed_13_0_426_inst_req_0;
      W_fetch_val_411_delayed_13_0_426_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_411_delayed_13_0_426_inst_req_1;
      W_fetch_val_411_delayed_13_0_426_inst_ack_1<= rack(0);
      W_fetch_val_411_delayed_13_0_426_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_411_delayed_13_0_426_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_411_delayed_13_0_428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_403_delayed_7_0_415_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_403_delayed_7_0_415_inst_req_0;
      W_fn_403_delayed_7_0_415_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_403_delayed_7_0_415_inst_req_1;
      W_fn_403_delayed_7_0_415_inst_ack_1<= rack(0);
      W_fn_403_delayed_7_0_415_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_403_delayed_7_0_415_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_403_delayed_7_0_417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_409_delayed_13_0_423_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_409_delayed_13_0_423_inst_req_0;
      W_fn_409_delayed_13_0_423_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_409_delayed_13_0_423_inst_req_1;
      W_fn_409_delayed_13_0_423_inst_ack_1<= rack(0);
      W_fn_409_delayed_13_0_423_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_409_delayed_13_0_423_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_409_delayed_13_0_425,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_344_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_344_final_reg_req_0;
      addr_of_344_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_344_final_reg_req_1;
      addr_of_344_final_reg_ack_1<= rack(0);
      addr_of_344_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_344_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_343_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_413_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_413_final_reg_req_0;
      addr_of_413_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_413_final_reg_req_1;
      addr_of_413_final_reg_ack_1<= rack(0);
      addr_of_413_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_413_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_412_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_349_368_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_349_368_buf_req_0;
      my_fetch_349_368_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_349_368_buf_req_1;
      my_fetch_349_368_buf_ack_1<= rack(0);
      my_fetch_349_368_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_349_368_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_349_368_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_434_369_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_434_369_buf_req_0;
      nfetch_val_434_369_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_434_369_buf_req_1;
      nfetch_val_434_369_buf_ack_1<= rack(0);
      nfetch_val_434_369_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_434_369_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_434_369_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_384_364_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_384_364_buf_req_0;
      nmycount_384_364_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_384_364_buf_req_1;
      nmycount_384_364_buf_ack_1<= rack(0);
      nmycount_384_364_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_384_364_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_384_364_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_365_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_365_buf_req_0;
      start_add_365_buf_ack_0<= wack(0);
      rreq(0) <= start_add_365_buf_req_1;
      start_add_365_buf_ack_1<= rack(0);
      start_add_365_buf : InterlockBuffer generic map ( -- 
        name => "start_add_365_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_365_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_337_inst
    process(pp_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := pp_buffer(0 downto 0);
      pingpong_338 <= tmp_var; -- 
    end process;
    -- interlock type_cast_389_inst
    process(LSHR_u64_u64_388_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_388_wire(15 downto 0);
      var_val_390 <= tmp_var; -- 
    end process;
    -- interlock type_cast_448_inst
    process(SUB_u64_u64_447_wire) -- 
      variable tmp_var : std_logic_vector(30 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 30 downto 0) := SUB_u64_u64_447_wire(30 downto 0);
      type_cast_448_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_343_index_1_rename
    process(R_sh_start_342_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_342_resized;
      ov(13 downto 0) := iv;
      R_sh_start_342_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_index_1_resize
    process(sh_start_334) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_334;
      ov := iv(13 downto 0);
      R_sh_start_342_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_343_root_address_inst
    process(array_obj_ref_343_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_343_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_343_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_index_1_rename
    process(LSHR_u64_u64_411_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_411_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_411_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_index_1_resize
    process(LSHR_u64_u64_411_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_411_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_411_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_412_root_address_inst
    process(array_obj_ref_412_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_412_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_412_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_348_addr_0
    process(ptr_deref_348_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_348_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_348_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_348_base_resize
    process(fetch_addr_345) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_345;
      ov := iv(13 downto 0);
      ptr_deref_348_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_348_gather_scatter
    process(ptr_deref_348_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_348_data_0;
      ov(63 downto 0) := iv;
      my_fetch_349 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_348_root_address_inst
    process(ptr_deref_348_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_348_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_348_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_421_addr_0
    process(ptr_deref_421_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_421_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_421_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_421_base_resize
    process(fetch_addr_414) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_414;
      ov := iv(13 downto 0);
      ptr_deref_421_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_421_gather_scatter
    process(ptr_deref_421_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_421_data_0;
      ov(63 downto 0) := iv;
      fv_422 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_421_root_address_inst
    process(ptr_deref_421_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_421_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_421_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_360_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_440_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_360_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_360_branch_req_0,
          ack0 => do_while_stmt_360_branch_ack_0,
          ack1 => do_while_stmt_360_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_383_inst
    process(mycount_362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_362, konst_382_wire_constant, tmp_var);
      nmycount_384 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_375_inst
    process(mycount_362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_362, konst_374_wire_constant, tmp_var);
      AND_u64_u64_375_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_402_inst
    process(nmycount_384) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_384, konst_401_wire_constant, tmp_var);
      AND_u64_u64_402_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : CONCAT_u1_u32_449_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pingpong_338 & type_cast_448_wire;
      CONCAT_u1_u32_449_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u32_449_inst_req_0;
      CONCAT_u1_u32_449_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u32_449_inst_req_1;
      CONCAT_u1_u32_449_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 31, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator EQ_u64_u1_353_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_352_wire_constant, tmp_var);
      first_fill_354 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_404_inst
    process(AND_u64_u64_402_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_402_wire, konst_403_wire_constant, tmp_var);
      fn_405 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_333_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_332_wire_constant, tmp_var);
      sh_start_334 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_388_inst
    process(fetch_val_366, my_num1_379) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_366, my_num1_379, tmp_var);
      LSHR_u64_u64_388_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_411_inst
    process(nmycount_384) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_384, konst_410_wire_constant, tmp_var);
      LSHR_u64_u64_411_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_378_inst
    process(SUB_u64_u64_376_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_376_wire, konst_377_wire_constant, tmp_var);
      my_num1_379 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_376_inst
    process(konst_372_wire_constant, AND_u64_u64_375_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_372_wire_constant, AND_u64_u64_375_wire, tmp_var);
      SUB_u64_u64_376_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_439_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_438_wire_constant, tmp_var);
      SUB_u64_u64_439_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_447_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_447_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_440_inst
    process(mycount_362, SUB_u64_u64_439_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_362, SUB_u64_u64_439_wire, tmp_var);
      ULT_u64_u1_440_wire <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_343_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_342_scaled;
      array_obj_ref_343_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_343_index_offset_req_0;
      array_obj_ref_343_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_343_index_offset_req_1;
      array_obj_ref_343_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : array_obj_ref_412_index_offset 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_411_scaled;
      array_obj_ref_412_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_412_index_offset_req_0;
      array_obj_ref_412_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_412_index_offset_req_1;
      array_obj_ref_412_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared load operator group (0) : ptr_deref_348_load_0 ptr_deref_421_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_348_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_421_load_0_req_0;
      ptr_deref_348_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_421_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_348_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_421_load_0_req_1;
      ptr_deref_348_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_421_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_403_delayed_7_0_417(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_348_word_address_0 & ptr_deref_421_word_address_0;
      ptr_deref_348_data_0 <= data_out(127 downto 64);
      ptr_deref_421_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_357_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_357_inst_req_0;
      RPIPE_input_done_pipe_357_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_357_inst_req_1;
      RPIPE_input_done_pipe_357_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_354(0);
      start_next_358 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_392_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_392_inst_req_0;
      WPIPE_kernel_pipe1_392_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_392_inst_req_1;
      WPIPE_kernel_pipe1_392_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not pingpong_338(0);
      data_in <= var_val_390;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_396_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_396_inst_req_0;
      WPIPE_kernel_pipe2_396_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_396_inst_req_1;
      WPIPE_kernel_pipe2_396_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= pingpong_338(0);
      data_in <= var_val_390;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_size_pipe_442_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_442_inst_req_0;
      WPIPE_size_pipe_442_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_442_inst_req_1;
      WPIPE_size_pipe_442_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u1_u32_449_wire;
      size_pipe_write_2_gI: SplitGuardInterface generic map(name => "size_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_318_inst_req_0 : boolean;
  signal WPIPE_timer_req_318_inst_ack_0 : boolean;
  signal WPIPE_timer_req_318_inst_req_1 : boolean;
  signal WPIPE_timer_req_318_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_323_inst_req_0 : boolean;
  signal RPIPE_timer_resp_323_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_323_inst_req_1 : boolean;
  signal RPIPE_timer_resp_323_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/req
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_sample_start_
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/rr
      -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => RPIPE_timer_resp_323_inst_req_0); -- 
    req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => WPIPE_timer_req_318_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_update_start_
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/ack
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/$entry
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/req
      -- 
    ack_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_318_inst_ack_0, ack => timer_CP_637_elements(1)); -- 
    req_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(1), ack => WPIPE_timer_req_318_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/ack
      -- 
    ack_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_318_inst_ack_1, ack => timer_CP_637_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_sample_completed_
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_update_start_
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/ra
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/$entry
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/cr
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_323_inst_ack_0, ack => timer_CP_637_elements(3)); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(3), ack => RPIPE_timer_resp_323_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_update_completed_
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/$exit
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_323_inst_ack_1, ack => timer_CP_637_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_321_to_assign_stmt_324/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_637_elements(2) & timer_CP_637_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_637_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_320_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_320_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_323_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_323_inst_req_0;
      RPIPE_timer_resp_323_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_323_inst_req_1;
      RPIPE_timer_resp_323_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_318_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_318_inst_req_0;
      WPIPE_timer_req_318_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_318_inst_req_1;
      WPIPE_timer_req_318_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_320_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4897_start: Boolean;
  signal timerDaemon_CP_4897_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2167_branch_req_0 : boolean;
  signal phi_stmt_2169_req_0 : boolean;
  signal phi_stmt_2169_req_1 : boolean;
  signal phi_stmt_2169_ack_0 : boolean;
  signal nCOUNTER_2182_2171_buf_req_0 : boolean;
  signal nCOUNTER_2182_2171_buf_ack_0 : boolean;
  signal nCOUNTER_2182_2171_buf_req_1 : boolean;
  signal nCOUNTER_2182_2171_buf_ack_1 : boolean;
  signal RPIPE_timer_req_2176_inst_req_0 : boolean;
  signal RPIPE_timer_req_2176_inst_ack_0 : boolean;
  signal RPIPE_timer_req_2176_inst_req_1 : boolean;
  signal RPIPE_timer_req_2176_inst_ack_1 : boolean;
  signal WPIPE_timer_resp_2184_inst_req_0 : boolean;
  signal WPIPE_timer_resp_2184_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_2184_inst_req_1 : boolean;
  signal WPIPE_timer_resp_2184_inst_ack_1 : boolean;
  signal do_while_stmt_2167_branch_ack_0 : boolean;
  signal do_while_stmt_2167_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4897_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4897_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4897_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4897_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4897: Block -- control-path 
    signal timerDaemon_CP_4897_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4897_elements(0) <= timerDaemon_CP_4897_start;
    timerDaemon_CP_4897_symbol <= timerDaemon_CP_4897_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2166/$entry
      -- CP-element group 0: 	 branch_block_stmt_2166/branch_block_stmt_2166__entry__
      -- CP-element group 0: 	 branch_block_stmt_2166/do_while_stmt_2167__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2166/$exit
      -- CP-element group 1: 	 branch_block_stmt_2166/branch_block_stmt_2166__exit__
      -- CP-element group 1: 	 branch_block_stmt_2166/do_while_stmt_2167__exit__
      -- 
    timerDaemon_CP_4897_elements(1) <= timerDaemon_CP_4897_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2166/do_while_stmt_2167/$entry
      -- CP-element group 2: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167__entry__
      -- 
    timerDaemon_CP_4897_elements(2) <= timerDaemon_CP_4897_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167__exit__
      -- 
    -- Element group timerDaemon_CP_4897_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_back
      -- 
    -- Element group timerDaemon_CP_4897_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2166/do_while_stmt_2167/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_taken/$entry
      -- 
    timerDaemon_CP_4897_elements(5) <= timerDaemon_CP_4897_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_body_done
      -- 
    timerDaemon_CP_4897_elements(6) <= timerDaemon_CP_4897_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4897_elements(7) <= timerDaemon_CP_4897_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4897_elements(8) <= timerDaemon_CP_4897_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2174_sample_start_
      -- 
    -- Element group timerDaemon_CP_4897_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/condition_evaluated
      -- 
    condition_evaluated_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(10), ack => do_while_stmt_2167_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(14) & timerDaemon_CP_4897_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(9) & timerDaemon_CP_4897_elements(15) & timerDaemon_CP_4897_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2174_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(35) & timerDaemon_CP_4897_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(32) & timerDaemon_CP_4897_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(18) & timerDaemon_CP_4897_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(9) & timerDaemon_CP_4897_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(9) & timerDaemon_CP_4897_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4897_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_4897_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_loopback_trigger
      -- 
    timerDaemon_CP_4897_elements(19) <= timerDaemon_CP_4897_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_loopback_sample_req_ps
      -- 
    phi_stmt_2169_loopback_sample_req_4936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2169_loopback_sample_req_4936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(20), ack => phi_stmt_2169_req_0); -- 
    -- Element group timerDaemon_CP_4897_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_entry_trigger
      -- 
    timerDaemon_CP_4897_elements(21) <= timerDaemon_CP_4897_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_entry_sample_req_ps
      -- 
    phi_stmt_2169_entry_sample_req_4939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2169_entry_sample_req_4939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(22), ack => phi_stmt_2169_req_1); -- 
    -- Element group timerDaemon_CP_4897_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2169_phi_mux_ack_ps
      -- 
    phi_stmt_2169_phi_mux_ack_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2169_ack_0, ack => timerDaemon_CP_4897_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Sample/req
      -- 
    req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(24), ack => nCOUNTER_2182_2171_buf_req_0); -- 
    -- Element group timerDaemon_CP_4897_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_update_start_
      -- CP-element group 25: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Update/req
      -- 
    req_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(25), ack => nCOUNTER_2182_2171_buf_req_1); -- 
    -- Element group timerDaemon_CP_4897_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Sample/ack
      -- 
    ack_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2182_2171_buf_ack_0, ack => timerDaemon_CP_4897_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/R_nCOUNTER_2171_Update/ack
      -- 
    ack_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2182_2171_buf_ack_1, ack => timerDaemon_CP_4897_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4897_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_update_start_
      -- 
    -- Element group timerDaemon_CP_4897_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_update_completed__ps
      -- 
    timerDaemon_CP_4897_elements(30) <= timerDaemon_CP_4897_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/type_cast_2173_update_completed_
      -- 
    -- Element group timerDaemon_CP_4897_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => timerDaemon_CP_4897_elements(29), ack => timerDaemon_CP_4897_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2174_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(9) & timerDaemon_CP_4897_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Sample/rr
      -- 
    rr_4982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(33), ack => RPIPE_timer_req_2176_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(11) & timerDaemon_CP_4897_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Update/cr
      -- 
    cr_4987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(34), ack => RPIPE_timer_req_2176_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(35) & timerDaemon_CP_4897_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Sample/ra
      -- 
    ra_4983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2176_inst_ack_0, ack => timerDaemon_CP_4897_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/phi_stmt_2174_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/RPIPE_timer_req_2176_Update/ca
      -- 
    ca_4988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2176_inst_ack_1, ack => timerDaemon_CP_4897_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Sample/req
      -- 
    req_4996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(37), ack => WPIPE_timer_resp_2184_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(18) & timerDaemon_CP_4897_elements(36) & timerDaemon_CP_4897_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Update/req
      -- 
    ack_4997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2184_inst_ack_0, ack => timerDaemon_CP_4897_elements(38)); -- 
    req_5001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4897_elements(38), ack => WPIPE_timer_resp_2184_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/WPIPE_timer_resp_2184_Update/ack
      -- 
    ack_5002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2184_inst_ack_1, ack => timerDaemon_CP_4897_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4897_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_4897_elements(9), ack => timerDaemon_CP_4897_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2166/do_while_stmt_2167/do_while_stmt_2167_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4897_elements(12) & timerDaemon_CP_4897_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4897_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_exit/ack
      -- 
    ack_5007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2167_branch_ack_0, ack => timerDaemon_CP_4897_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_2166/do_while_stmt_2167/loop_taken/ack
      -- 
    ack_5011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2167_branch_ack_1, ack => timerDaemon_CP_4897_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2166/do_while_stmt_2167/$exit
      -- 
    timerDaemon_CP_4897_elements(44) <= timerDaemon_CP_4897_elements(3);
    timerDaemon_do_while_stmt_2167_terminator_5012: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2167_terminator_5012", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_4897_elements(6),loop_continue => timerDaemon_CP_4897_elements(43),loop_terminate => timerDaemon_CP_4897_elements(42),loop_back => timerDaemon_CP_4897_elements(4),loop_exit => timerDaemon_CP_4897_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2169_phi_seq_4970_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4897_elements(19);
      timerDaemon_CP_4897_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4897_elements(26);
      timerDaemon_CP_4897_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4897_elements(27);
      timerDaemon_CP_4897_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4897_elements(21);
      timerDaemon_CP_4897_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4897_elements(28);
      timerDaemon_CP_4897_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4897_elements(30);
      timerDaemon_CP_4897_elements(22) <= phi_mux_reqs(1);
      phi_stmt_2169_phi_seq_4970 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2169_phi_seq_4970") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4897_elements(11), 
          phi_sample_ack => timerDaemon_CP_4897_elements(17), 
          phi_update_req => timerDaemon_CP_4897_elements(13), 
          phi_update_ack => timerDaemon_CP_4897_elements(18), 
          phi_mux_ack => timerDaemon_CP_4897_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4922_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4897_elements(7);
        preds(1)  <= timerDaemon_CP_4897_elements(8);
        entry_tmerge_4922 : transition_merge -- 
          generic map(name => " entry_tmerge_4922")
          port map (preds => preds, symbol_out => timerDaemon_CP_4897_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2169 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_2176_wire : std_logic_vector(0 downto 0);
    signal konst_2180_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2188_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_2182 : std_logic_vector(63 downto 0);
    signal nCOUNTER_2182_2171_buffered : std_logic_vector(63 downto 0);
    signal req_2174 : std_logic_vector(0 downto 0);
    signal type_cast_2173_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_2180_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2188_wire_constant <= "1";
    type_cast_2173_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2169: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nCOUNTER_2182_2171_buffered & type_cast_2173_wire_constant;
      req <= phi_stmt_2169_req_0 & phi_stmt_2169_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2169",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2169_ack_0,
          idata => idata,
          odata => COUNTER_2169,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2169
    nCOUNTER_2182_2171_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_2182_2171_buf_req_0;
      nCOUNTER_2182_2171_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_2182_2171_buf_req_1;
      nCOUNTER_2182_2171_buf_ack_1<= rack(0);
      nCOUNTER_2182_2171_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_2182_2171_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_2182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_2182_2171_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2174
    process(RPIPE_timer_req_2176_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_2176_wire(0 downto 0);
      req_2174 <= tmp_var; -- 
    end process;
    do_while_stmt_2167_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2188_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2167_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2167_branch_req_0,
          ack0 => do_while_stmt_2167_branch_ack_0,
          ack1 => do_while_stmt_2167_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_2181_inst
    process(COUNTER_2169) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2169, konst_2180_wire_constant, tmp_var);
      nCOUNTER_2182 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_2176_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_2176_inst_req_0;
      RPIPE_timer_req_2176_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_2176_inst_req_1;
      RPIPE_timer_req_2176_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_2176_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_2184_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_2184_inst_req_0;
      WPIPE_timer_resp_2184_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_2184_inst_req_1;
      WPIPE_timer_resp_2184_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_2174(0);
      data_in <= COUNTER_2169;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(135 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      pp : in  std_logic_vector(7 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_pp :  std_logic_vector(7 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(135 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(135 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(135 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(135 downto 72);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(71 downto 8);
  loadKernelChannel_pp <= loadKernelChannel_in_args(7 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 136,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      pp => loadKernelChannel_pp,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(1 downto 1),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(1 downto 1),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
