-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_T;
architecture fill_T_arch of fill_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_T_CP_0_start: Boolean;
  signal fill_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_38_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_38_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_38_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_38_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_40_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_40_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_40_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_40_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_43_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_43_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_43_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_43_inst_ack_1 : boolean;
  signal CONCAT_u240_u256_56_inst_req_0 : boolean;
  signal CONCAT_u240_u256_56_inst_ack_0 : boolean;
  signal CONCAT_u240_u256_56_inst_req_1 : boolean;
  signal CONCAT_u240_u256_56_inst_ack_1 : boolean;
  signal if_stmt_58_branch_req_0 : boolean;
  signal if_stmt_58_branch_ack_1 : boolean;
  signal if_stmt_58_branch_ack_0 : boolean;
  signal phi_stmt_17_req_1 : boolean;
  signal phi_stmt_23_req_1 : boolean;
  signal nmycount_33_19_buf_req_0 : boolean;
  signal nmycount_33_19_buf_ack_0 : boolean;
  signal nmycount_33_19_buf_req_1 : boolean;
  signal nmycount_33_19_buf_ack_1 : boolean;
  signal phi_stmt_17_req_0 : boolean;
  signal ninput_word_57_25_buf_req_0 : boolean;
  signal ninput_word_57_25_buf_ack_0 : boolean;
  signal ninput_word_57_25_buf_req_1 : boolean;
  signal ninput_word_57_25_buf_ack_1 : boolean;
  signal phi_stmt_23_req_0 : boolean;
  signal phi_stmt_17_ack_0 : boolean;
  signal phi_stmt_23_ack_0 : boolean;
  signal array_obj_ref_71_index_offset_req_0 : boolean;
  signal array_obj_ref_71_index_offset_ack_0 : boolean;
  signal array_obj_ref_71_index_offset_req_1 : boolean;
  signal array_obj_ref_71_index_offset_ack_1 : boolean;
  signal addr_of_72_final_reg_req_0 : boolean;
  signal addr_of_72_final_reg_ack_0 : boolean;
  signal addr_of_72_final_reg_req_1 : boolean;
  signal addr_of_72_final_reg_ack_1 : boolean;
  signal ptr_deref_75_store_0_req_0 : boolean;
  signal ptr_deref_75_store_0_ack_0 : boolean;
  signal ptr_deref_75_store_0_req_1 : boolean;
  signal ptr_deref_75_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_T_CP_0: Block -- control-path 
    signal fill_T_CP_0_elements: BooleanArray(37 downto 0);
    -- 
  begin -- 
    fill_T_CP_0_elements(0) <= fill_T_CP_0_start;
    fill_T_CP_0_symbol <= fill_T_CP_0_elements(37);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	16 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_15/$entry
      -- CP-element group 0: 	 branch_block_stmt_15/branch_block_stmt_15__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	30 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1: 	12 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_15/merge_stmt_16__exit__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57__entry__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_update_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Update/cr
      -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => RPIPE_maxpool_input_pipe_35_inst_req_0); -- 
    cr_85_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_85_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u240_u256_56_inst_req_1); -- 
    fill_T_CP_0_elements(1) <= fill_T_CP_0_elements(30);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_update_start_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Sample/$exit
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_35_inst_ack_0, ack => fill_T_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(2), ack => RPIPE_maxpool_input_pipe_35_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_35_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Sample/req
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_35_inst_ack_1, ack => fill_T_CP_0_elements(3)); -- 
    rr_38_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_38_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => RPIPE_maxpool_input_pipe_38_inst_req_0); -- 
    req_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => WPIPE_maxpool_output_pipe_40_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_update_start_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Update/cr
      -- 
    ra_39_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_38_inst_ack_0, ack => fill_T_CP_0_elements(4)); -- 
    cr_43_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_43_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(4), ack => RPIPE_maxpool_input_pipe_38_inst_req_1); -- 
    -- CP-element group 5:  fork  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/RPIPE_maxpool_input_pipe_38_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Sample/rr
      -- 
    ca_44_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_38_inst_ack_1, ack => fill_T_CP_0_elements(5)); -- 
    rr_80_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_80_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(5), ack => CONCAT_u240_u256_56_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_update_start_
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Sample/ack
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Update/req
      -- 
    ack_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_40_inst_ack_0, ack => fill_T_CP_0_elements(6)); -- 
    req_57_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_57_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(6), ack => WPIPE_maxpool_output_pipe_40_inst_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_40_Update/ack
      -- 
    ack_58_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_40_inst_ack_1, ack => fill_T_CP_0_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Sample/req
      -- 
    req_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(8), ack => WPIPE_maxpool_output_pipe_43_inst_req_0); -- 
    fill_T_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "fill_T_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(7) & fill_T_CP_0_elements(5);
      gj_fill_T_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_update_start_
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Update/req
      -- 
    ack_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_43_inst_ack_0, ack => fill_T_CP_0_elements(9)); -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(9), ack => WPIPE_maxpool_output_pipe_43_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/WPIPE_maxpool_output_pipe_43_Update/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_43_inst_ack_1, ack => fill_T_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Sample/ra
      -- 
    ra_81_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_56_inst_ack_0, ack => fill_T_CP_0_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	1 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/CONCAT_u240_u256_56_Update/ca
      -- 
    ca_86_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_56_inst_ack_1, ack => fill_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  branch  join  transition  place  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (24) 
      -- CP-element group 13: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57__exit__
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58__entry__
      -- CP-element group 13: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_57/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/ULT_u4_u1_61_inputs/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/ULT_u4_u1_61_inputs/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Update/cr
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/ULT_u4_u1_61/SplitProtocol/Update/ca
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_15/ULT_u4_u1_61_place
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_15/if_stmt_58_else_link/$entry
      -- 
    branch_req_113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(13), ack => if_stmt_58_branch_req_0); -- 
    fill_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(10) & fill_T_CP_0_elements(12);
      gj_fill_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	23 
    -- CP-element group 14: 	24 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14:  members (18) 
      -- CP-element group 14: 	 branch_block_stmt_15/if_stmt_58_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_15/if_stmt_58_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_15/loopback
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/req
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/req
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/req
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/req
      -- 
    if_choice_transition_118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_58_branch_ack_1, ack => fill_T_CP_0_elements(14)); -- 
    req_162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => nmycount_33_19_buf_req_0); -- 
    req_167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => nmycount_33_19_buf_req_1); -- 
    req_182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => ninput_word_57_25_buf_req_0); -- 
    req_187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => ninput_word_57_25_buf_req_1); -- 
    -- CP-element group 15:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	36 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	34 
    -- CP-element group 15:  members (30) 
      -- CP-element group 15: 	 branch_block_stmt_15/$exit
      -- CP-element group 15: 	 branch_block_stmt_15/branch_block_stmt_15__exit__
      -- CP-element group 15: 	 branch_block_stmt_15/if_stmt_58__exit__
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_scale_1/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_scale_1/$exit
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_scale_1/scale_rename_req
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_scale_1/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_15/if_stmt_58_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_15/if_stmt_58_else_link/else_choice_transition
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_update_start_
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_resized_1
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_scaled_1
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_computed_1
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_resize_1/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_resize_1/$exit
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_resize_1/index_resize_req
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_index_resize_1/index_resize_ack
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_update_start
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Sample/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Sample/req
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Update/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Update/req
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_complete/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_complete/req
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_update_start_
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_58_branch_ack_0, ack => fill_T_CP_0_elements(15)); -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(15), ack => array_obj_ref_71_index_offset_req_0); -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(15), ack => array_obj_ref_71_index_offset_req_1); -- 
    req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(15), ack => addr_of_72_final_reg_req_1); -- 
    cr_293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(15), ack => ptr_deref_75_store_0_req_1); -- 
    -- CP-element group 16:  fork  transition  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$entry
      -- CP-element group 16: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$entry
      -- CP-element group 16: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 16: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$entry
      -- CP-element group 16: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- 
    fill_T_CP_0_elements(16) <= fill_T_CP_0_elements(0);
    -- CP-element group 17:  transition  output  delay-element  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$exit
      -- CP-element group 17: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 17: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/type_cast_22_konst_delay_trans
      -- CP-element group 17: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(17), ack => phi_stmt_17_req_1); -- 
    -- Element group fill_T_CP_0_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(16), ack => fill_T_CP_0_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  transition  output  delay-element  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/type_cast_27_konst_delay_trans
      -- CP-element group 18: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(18), ack => phi_stmt_23_req_1); -- 
    -- Element group fill_T_CP_0_elements(18) is a control-delay.
    cp_element_18_delay: control_delay_element  generic map(name => " 18_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(16), ack => fill_T_CP_0_elements(18), clk => clk, reset =>reset);
    -- CP-element group 19:  join  transition  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	27 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$exit
      -- 
    fill_T_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(18) & fill_T_CP_0_elements(17);
      gj_fill_T_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/ack
      -- 
    ack_163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_19_buf_ack_0, ack => fill_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/ack
      -- 
    ack_168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_19_buf_ack_1, ack => fill_T_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	26 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$exit
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$exit
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(22), ack => phi_stmt_17_req_0); -- 
    fill_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(20) & fill_T_CP_0_elements(21);
      gj_fill_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	14 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/ack
      -- 
    ack_183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_57_25_buf_ack_0, ack => fill_T_CP_0_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	14 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/ack
      -- 
    ack_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_57_25_buf_ack_1, ack => fill_T_CP_0_elements(24)); -- 
    -- CP-element group 25:  join  transition  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$exit
      -- CP-element group 25: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 25: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$exit
      -- CP-element group 25: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(25), ack => phi_stmt_23_req_0); -- 
    fill_T_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(23) & fill_T_CP_0_elements(24);
      gj_fill_T_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: 	22 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_15/loopback_PhiReq/$exit
      -- 
    fill_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(25) & fill_T_CP_0_elements(22);
      gj_fill_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  merge  fork  transition  place  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_15/merge_stmt_16_PhiReqMerge
      -- CP-element group 27: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$entry
      -- 
    fill_T_CP_0_elements(27) <= OrReduce(fill_T_CP_0_elements(19) & fill_T_CP_0_elements(26));
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_17_ack
      -- 
    phi_stmt_17_ack_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_17_ack_0, ack => fill_T_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_23_ack
      -- 
    phi_stmt_23_ack_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_23_ack_0, ack => fill_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  transition  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	1 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$exit
      -- 
    fill_T_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(28) & fill_T_CP_0_elements(29);
      gj_fill_T_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	37 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_sample_complete
      -- CP-element group 31: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_offset_ack_0, ack => fill_T_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (11) 
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_sample_start_
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_root_address_calculated
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_offset_calculated
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Update/$exit
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_final_index_sum_regn_Update/ack
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_base_plus_offset/$entry
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_base_plus_offset/$exit
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_base_plus_offset/sum_rename_req
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/array_obj_ref_71_base_plus_offset/sum_rename_ack
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_request/$entry
      -- CP-element group 32: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_request/req
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_71_index_offset_ack_1, ack => fill_T_CP_0_elements(32)); -- 
    req_238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(32), ack => addr_of_72_final_reg_req_0); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_sample_completed_
      -- CP-element group 33: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_request/$exit
      -- CP-element group 33: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_request/ack
      -- 
    ack_239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_72_final_reg_ack_0, ack => fill_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	15 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_update_completed_
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_complete/$exit
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/addr_of_72_complete/ack
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_sample_start_
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_address_calculated
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_word_address_calculated
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_root_address_calculated
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_address_resized
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_addr_resize/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_addr_resize/$exit
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_addr_resize/base_resize_req
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_addr_resize/base_resize_ack
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_plus_offset/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_plus_offset/$exit
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_plus_offset/sum_rename_req
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_base_plus_offset/sum_rename_ack
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_word_addrgen/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_word_addrgen/$exit
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_word_addrgen/root_register_req
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_word_addrgen/root_register_ack
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/ptr_deref_75_Split/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/ptr_deref_75_Split/$exit
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/ptr_deref_75_Split/split_req
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/ptr_deref_75_Split/split_ack
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/word_0/$entry
      -- CP-element group 34: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/word_0/rr
      -- 
    ack_244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_72_final_reg_ack_1, ack => fill_T_CP_0_elements(34)); -- 
    rr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(34), ack => ptr_deref_75_store_0_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (5) 
      -- CP-element group 35: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_sample_completed_
      -- CP-element group 35: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/$exit
      -- CP-element group 35: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/$exit
      -- CP-element group 35: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/word_0/$exit
      -- CP-element group 35: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Sample/word_access_start/word_0/ra
      -- 
    ra_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_75_store_0_ack_0, ack => fill_T_CP_0_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	15 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_update_completed_
      -- CP-element group 36: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/$exit
      -- CP-element group 36: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/$exit
      -- CP-element group 36: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/word_0/$exit
      -- CP-element group 36: 	 assign_stmt_73_to_assign_stmt_77/ptr_deref_75_Update/word_access_complete/word_0/ca
      -- 
    ca_294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_75_store_0_ack_1, ack => fill_T_CP_0_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	31 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 $exit
      -- CP-element group 37: 	 assign_stmt_73_to_assign_stmt_77/$exit
      -- 
    fill_T_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(36) & fill_T_CP_0_elements(31);
      gj_fill_T_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(37), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_addr_70_resized : std_logic_vector(13 downto 0);
    signal R_addr_70_scaled : std_logic_vector(13 downto 0);
    signal ULT_u4_u1_61_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_71_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_71_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_71_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_71_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_71_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_71_root_address : std_logic_vector(13 downto 0);
    signal input_word_23 : std_logic_vector(255 downto 0);
    signal konst_31_wire_constant : std_logic_vector(3 downto 0);
    signal konst_60_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_17 : std_logic_vector(3 downto 0);
    signal ninput_word_57 : std_logic_vector(255 downto 0);
    signal ninput_word_57_25_buffered : std_logic_vector(255 downto 0);
    signal nmycount_33 : std_logic_vector(3 downto 0);
    signal nmycount_33_19_buffered : std_logic_vector(3 downto 0);
    signal ptr_73 : std_logic_vector(31 downto 0);
    signal ptr_deref_75_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_75_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_75_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_75_wire : std_logic_vector(255 downto 0);
    signal ptr_deref_75_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_75_word_offset_0 : std_logic_vector(13 downto 0);
    signal slice_54_wire : std_logic_vector(239 downto 0);
    signal type_cast_22_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_27_wire_constant : std_logic_vector(255 downto 0);
    signal val1_36 : std_logic_vector(7 downto 0);
    signal val2_39 : std_logic_vector(7 downto 0);
    signal val_50 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_71_constant_part_of_offset <= "00000000000000";
    array_obj_ref_71_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_71_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_71_resized_base_address <= "00000000000000";
    konst_31_wire_constant <= "0001";
    konst_60_wire_constant <= "1111";
    ptr_deref_75_word_offset_0 <= "00000000000000";
    type_cast_22_wire_constant <= "0000";
    type_cast_27_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_17: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_33_19_buffered & type_cast_22_wire_constant;
      req <= phi_stmt_17_req_0 & phi_stmt_17_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_17",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_17_ack_0,
          idata => idata,
          odata => mycount_17,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_17
    phi_stmt_23: Block -- phi operator 
      signal idata: std_logic_vector(511 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ninput_word_57_25_buffered & type_cast_27_wire_constant;
      req <= phi_stmt_23_req_0 & phi_stmt_23_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_23",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 256) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_23_ack_0,
          idata => idata,
          odata => input_word_23,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_23
    -- flow-through slice operator slice_54_inst
    slice_54_wire <= input_word_23(239 downto 0);
    addr_of_72_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_72_final_reg_req_0;
      addr_of_72_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_72_final_reg_req_1;
      addr_of_72_final_reg_ack_1<= rack(0);
      addr_of_72_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_72_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_71_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_73,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ninput_word_57_25_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_57_25_buf_req_0;
      ninput_word_57_25_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_57_25_buf_req_1;
      ninput_word_57_25_buf_ack_1<= rack(0);
      ninput_word_57_25_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_57_25_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 256,
        out_data_width => 256,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_57,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_57_25_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_33_19_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_33_19_buf_req_0;
      nmycount_33_19_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_33_19_buf_req_1;
      nmycount_33_19_buf_ack_1<= rack(0);
      nmycount_33_19_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_33_19_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_33,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_33_19_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_71_index_1_rename
    process(R_addr_70_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_70_resized;
      ov(13 downto 0) := iv;
      R_addr_70_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_70_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_71_root_address_inst
    process(array_obj_ref_71_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_71_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_71_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_75_addr_0
    process(ptr_deref_75_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_75_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_75_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_75_base_resize
    process(ptr_73) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_73;
      ov := iv(13 downto 0);
      ptr_deref_75_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_75_gather_scatter
    process(ninput_word_57) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_57;
      ov(255 downto 0) := iv;
      ptr_deref_75_data_0 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_75_root_address_inst
    process(ptr_deref_75_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_75_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_75_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_58_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_61_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_58_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_58_branch_req_0,
          ack0 => if_stmt_58_branch_ack_0,
          ack1 => if_stmt_58_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u4_u4_32_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_17, konst_31_wire_constant, tmp_var);
      nmycount_33 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u240_u256_56_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_54_wire & val_50;
      ninput_word_57 <= data_out(255 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u240_u256_56_inst_req_0;
      CONCAT_u240_u256_56_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u240_u256_56_inst_req_1;
      CONCAT_u240_u256_56_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 240,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 256,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator CONCAT_u8_u16_49_inst
    process(val1_36, val2_39) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(val1_36, val2_39, tmp_var);
      val_50 <= tmp_var; --
    end process;
    -- binary operator ULT_u4_u1_61_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_17, konst_60_wire_constant, tmp_var);
      ULT_u4_u1_61_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_71_index_offset 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_70_scaled;
      array_obj_ref_71_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_71_index_offset_req_0;
      array_obj_ref_71_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_71_index_offset_req_1;
      array_obj_ref_71_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared store operator group (0) : ptr_deref_75_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_75_store_0_req_0;
      ptr_deref_75_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_75_store_0_req_1;
      ptr_deref_75_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_75_word_address_0;
      data_in <= ptr_deref_75_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 256,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(255 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_35_inst RPIPE_maxpool_input_pipe_38_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_35_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_38_inst_req_0;
      RPIPE_maxpool_input_pipe_35_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_38_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_35_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_38_inst_req_1;
      RPIPE_maxpool_input_pipe_35_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_38_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      val1_36 <= data_out(15 downto 8);
      val2_39 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_40_inst WPIPE_maxpool_output_pipe_43_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_40_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_43_inst_req_0;
      WPIPE_maxpool_output_pipe_40_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_43_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_40_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_43_inst_req_1;
      WPIPE_maxpool_output_pipe_40_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_43_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= val1_36 & val2_39;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    fill_T_call_reqs : out  std_logic_vector(0 downto 0);
    fill_T_call_acks : in   std_logic_vector(0 downto 0);
    fill_T_call_data : out  std_logic_vector(63 downto 0);
    fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_T_return_reqs : out  std_logic_vector(0 downto 0);
    fill_T_return_acks : in   std_logic_vector(0 downto 0);
    fill_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(159 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool3D;
architecture maxPool3D_arch of maxPool3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal maxPool3D_CP_2672_start: Boolean;
  signal maxPool3D_CP_2672_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_1672_inst_req_1 : boolean;
  signal type_cast_1667_inst_req_1 : boolean;
  signal type_cast_1363_inst_req_0 : boolean;
  signal type_cast_1622_inst_ack_1 : boolean;
  signal type_cast_1363_inst_req_1 : boolean;
  signal type_cast_1363_inst_ack_0 : boolean;
  signal type_cast_1672_inst_ack_1 : boolean;
  signal type_cast_1681_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1346_inst_req_0 : boolean;
  signal W_colx_x1_1760_delayed_1_0_1770_inst_req_0 : boolean;
  signal type_cast_1363_inst_ack_1 : boolean;
  signal type_cast_1667_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_req_1 : boolean;
  signal type_cast_1667_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1396_inst_ack_1 : boolean;
  signal phi_stmt_1659_ack_0 : boolean;
  signal type_cast_1350_inst_ack_1 : boolean;
  signal W_rowx_x1_1781_delayed_2_0_1794_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_ack_1 : boolean;
  signal type_cast_1400_inst_req_0 : boolean;
  signal type_cast_1400_inst_ack_0 : boolean;
  signal type_cast_1350_inst_req_1 : boolean;
  signal type_cast_1768_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1396_inst_req_1 : boolean;
  signal type_cast_1350_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_ack_0 : boolean;
  signal type_cast_1350_inst_req_0 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal type_cast_1672_inst_req_0 : boolean;
  signal type_cast_1375_inst_ack_1 : boolean;
  signal type_cast_1672_inst_ack_0 : boolean;
  signal type_cast_1375_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_1 : boolean;
  signal type_cast_1768_inst_ack_1 : boolean;
  signal type_cast_1400_inst_ack_1 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal type_cast_1375_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_0 : boolean;
  signal type_cast_1400_inst_req_1 : boolean;
  signal type_cast_1375_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_0 : boolean;
  signal W_rowx_x1_1781_delayed_2_0_1794_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1396_inst_ack_0 : boolean;
  signal phi_stmt_1659_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_ack_0 : boolean;
  signal type_cast_1622_inst_req_1 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1346_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1371_inst_req_0 : boolean;
  signal W_rowx_x1_1781_delayed_2_0_1794_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1346_inst_req_1 : boolean;
  signal type_cast_1768_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1396_inst_req_0 : boolean;
  signal do_while_stmt_1657_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1346_inst_ack_0 : boolean;
  signal phi_stmt_1659_req_1 : boolean;
  signal phi_stmt_1664_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1409_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1409_inst_ack_0 : boolean;
  signal if_stmt_1820_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1409_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1409_inst_ack_1 : boolean;
  signal type_cast_1681_inst_req_1 : boolean;
  signal type_cast_1413_inst_req_0 : boolean;
  signal type_cast_1413_inst_ack_0 : boolean;
  signal type_cast_1413_inst_req_1 : boolean;
  signal type_cast_1413_inst_ack_1 : boolean;
  signal call_stmt_1833_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1421_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1421_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1421_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1421_inst_ack_1 : boolean;
  signal type_cast_1681_inst_ack_0 : boolean;
  signal type_cast_1662_inst_ack_1 : boolean;
  signal type_cast_1681_inst_req_0 : boolean;
  signal type_cast_1662_inst_req_1 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal call_stmt_1833_call_req_1 : boolean;
  signal call_stmt_1754_call_ack_1 : boolean;
  signal call_stmt_1754_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1434_inst_ack_1 : boolean;
  signal type_cast_1438_inst_req_0 : boolean;
  signal phi_stmt_1669_ack_0 : boolean;
  signal type_cast_1438_inst_ack_0 : boolean;
  signal type_cast_1792_inst_ack_1 : boolean;
  signal type_cast_1438_inst_req_1 : boolean;
  signal type_cast_1438_inst_ack_1 : boolean;
  signal type_cast_1837_inst_ack_0 : boolean;
  signal call_stmt_1754_call_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1446_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1446_inst_ack_0 : boolean;
  signal type_cast_1829_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1446_inst_req_1 : boolean;
  signal phi_stmt_1669_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1446_inst_ack_1 : boolean;
  signal type_cast_1662_inst_ack_0 : boolean;
  signal type_cast_1662_inst_req_0 : boolean;
  signal type_cast_1792_inst_req_1 : boolean;
  signal type_cast_1450_inst_req_0 : boolean;
  signal type_cast_1450_inst_ack_0 : boolean;
  signal type_cast_1450_inst_req_1 : boolean;
  signal type_cast_1450_inst_ack_1 : boolean;
  signal type_cast_1837_inst_req_0 : boolean;
  signal call_stmt_1754_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_req_0 : boolean;
  signal phi_stmt_1669_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_ack_0 : boolean;
  signal type_cast_1829_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1459_inst_ack_1 : boolean;
  signal type_cast_1677_inst_ack_1 : boolean;
  signal type_cast_1677_inst_req_1 : boolean;
  signal type_cast_1463_inst_req_0 : boolean;
  signal type_cast_1463_inst_ack_0 : boolean;
  signal type_cast_1792_inst_ack_0 : boolean;
  signal type_cast_1463_inst_req_1 : boolean;
  signal type_cast_1463_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1471_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1471_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1471_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1471_inst_ack_1 : boolean;
  signal type_cast_1677_inst_ack_0 : boolean;
  signal type_cast_1792_inst_req_0 : boolean;
  signal type_cast_1475_inst_req_0 : boolean;
  signal type_cast_1475_inst_ack_0 : boolean;
  signal type_cast_1475_inst_req_1 : boolean;
  signal type_cast_1475_inst_ack_1 : boolean;
  signal type_cast_1677_inst_req_0 : boolean;
  signal type_cast_1685_inst_ack_1 : boolean;
  signal type_cast_1685_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1484_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1484_inst_ack_0 : boolean;
  signal type_cast_1829_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1484_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1484_inst_ack_1 : boolean;
  signal do_while_stmt_1657_branch_ack_1 : boolean;
  signal type_cast_1488_inst_req_0 : boolean;
  signal type_cast_1488_inst_ack_0 : boolean;
  signal type_cast_1488_inst_req_1 : boolean;
  signal type_cast_1488_inst_ack_1 : boolean;
  signal call_stmt_1833_call_ack_0 : boolean;
  signal if_stmt_1820_branch_ack_0 : boolean;
  signal type_cast_1498_inst_req_0 : boolean;
  signal type_cast_1498_inst_ack_0 : boolean;
  signal type_cast_1498_inst_req_1 : boolean;
  signal type_cast_1498_inst_ack_1 : boolean;
  signal call_stmt_1833_call_req_0 : boolean;
  signal type_cast_1626_inst_ack_1 : boolean;
  signal if_stmt_1516_branch_req_0 : boolean;
  signal do_while_stmt_1657_branch_ack_0 : boolean;
  signal type_cast_1626_inst_req_1 : boolean;
  signal if_stmt_1516_branch_ack_1 : boolean;
  signal if_stmt_1516_branch_ack_0 : boolean;
  signal type_cast_1829_inst_req_0 : boolean;
  signal type_cast_1768_inst_ack_0 : boolean;
  signal W_colx_x1_1760_delayed_1_0_1770_inst_ack_1 : boolean;
  signal type_cast_1553_inst_req_0 : boolean;
  signal type_cast_1553_inst_ack_0 : boolean;
  signal phi_stmt_1664_ack_0 : boolean;
  signal W_colx_x1_1760_delayed_1_0_1770_inst_req_1 : boolean;
  signal type_cast_1553_inst_req_1 : boolean;
  signal type_cast_1553_inst_ack_1 : boolean;
  signal if_stmt_1820_branch_ack_1 : boolean;
  signal type_cast_1685_inst_ack_0 : boolean;
  signal W_colx_x1_1760_delayed_1_0_1770_inst_ack_0 : boolean;
  signal call_stmt_1579_call_req_0 : boolean;
  signal call_stmt_1579_call_ack_0 : boolean;
  signal call_stmt_1579_call_req_1 : boolean;
  signal call_stmt_1579_call_ack_1 : boolean;
  signal type_cast_1837_inst_req_1 : boolean;
  signal type_cast_1685_inst_req_0 : boolean;
  signal type_cast_1626_inst_ack_0 : boolean;
  signal if_stmt_1591_branch_req_0 : boolean;
  signal type_cast_1626_inst_req_0 : boolean;
  signal phi_stmt_1664_req_1 : boolean;
  signal if_stmt_1591_branch_ack_1 : boolean;
  signal if_stmt_1591_branch_ack_0 : boolean;
  signal W_rowx_x1_1781_delayed_2_0_1794_inst_ack_1 : boolean;
  signal call_stmt_1614_call_req_0 : boolean;
  signal type_cast_1667_inst_ack_1 : boolean;
  signal call_stmt_1614_call_ack_0 : boolean;
  signal call_stmt_1614_call_req_1 : boolean;
  signal call_stmt_1614_call_ack_1 : boolean;
  signal type_cast_1618_inst_req_0 : boolean;
  signal type_cast_1618_inst_ack_0 : boolean;
  signal type_cast_1618_inst_req_1 : boolean;
  signal type_cast_1618_inst_ack_1 : boolean;
  signal type_cast_1622_inst_req_0 : boolean;
  signal type_cast_1622_inst_ack_0 : boolean;
  signal type_cast_1837_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1844_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1844_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1844_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1844_inst_ack_1 : boolean;
  signal type_cast_1850_inst_req_0 : boolean;
  signal type_cast_1850_inst_ack_0 : boolean;
  signal type_cast_1850_inst_req_1 : boolean;
  signal type_cast_1850_inst_ack_1 : boolean;
  signal type_cast_1854_inst_req_0 : boolean;
  signal type_cast_1854_inst_ack_0 : boolean;
  signal type_cast_1854_inst_req_1 : boolean;
  signal type_cast_1854_inst_ack_1 : boolean;
  signal call_stmt_1867_call_req_0 : boolean;
  signal call_stmt_1867_call_ack_0 : boolean;
  signal call_stmt_1867_call_req_1 : boolean;
  signal call_stmt_1867_call_ack_1 : boolean;
  signal phi_stmt_1570_req_0 : boolean;
  signal type_cast_1576_inst_req_0 : boolean;
  signal type_cast_1576_inst_ack_0 : boolean;
  signal type_cast_1576_inst_req_1 : boolean;
  signal type_cast_1576_inst_ack_1 : boolean;
  signal phi_stmt_1570_req_1 : boolean;
  signal phi_stmt_1570_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool3D_CP_2672_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2672_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool3D_CP_2672_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2672_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool3D_CP_2672: Block -- control-path 
    signal maxPool3D_CP_2672_elements: BooleanArray(204 downto 0);
    -- 
  begin -- 
    maxPool3D_CP_2672_elements(0) <= maxPool3D_CP_2672_start;
    maxPool3D_CP_2672_symbol <= maxPool3D_CP_2672_elements(197);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0:  members (44) 
      -- CP-element group 0: 	 branch_block_stmt_1344/branch_block_stmt_1344__entry__
      -- CP-element group 0: 	 branch_block_stmt_1344/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494__entry__
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Update/cr
      -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1363_inst_req_1); -- 
    rr_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => RPIPE_maxpool_input_pipe_1346_inst_req_0); -- 
    cr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1350_inst_req_1); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1375_inst_req_1); -- 
    cr_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1388_inst_req_1); -- 
    cr_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1400_inst_req_1); -- 
    cr_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1413_inst_req_1); -- 
    cr_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1425_inst_req_1); -- 
    cr_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1438_inst_req_1); -- 
    cr_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1450_inst_req_1); -- 
    cr_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1463_inst_req_1); -- 
    cr_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1475_inst_req_1); -- 
    cr_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(0), ack => type_cast_1488_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	180 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	181 
    -- CP-element group 1: 	182 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820__entry__
      -- CP-element group 1: 	 branch_block_stmt_1344/do_while_stmt_1657__exit__
      -- CP-element group 1: 	 branch_block_stmt_1344/R_whilex_xbody_whilex_xend_taken_1821_place
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1344/if_stmt_1820_else_link/$entry
      -- 
    branch_req_3496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(1), ack => if_stmt_1820_branch_req_0); -- 
    maxPool3D_CP_2672_elements(1) <= maxPool3D_CP_2672_elements(180);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Sample/ra
      -- 
    ra_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1346_inst_ack_0, ack => maxPool3D_CP_2672_elements(2)); -- 
    cr_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(2), ack => RPIPE_maxpool_input_pipe_1346_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1346_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_sample_start_
      -- 
    ca_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1346_inst_ack_1, ack => maxPool3D_CP_2672_elements(3)); -- 
    rr_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(3), ack => type_cast_1350_inst_req_0); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(3), ack => RPIPE_maxpool_input_pipe_1359_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_sample_completed_
      -- 
    ra_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1350_inst_ack_0, ack => maxPool3D_CP_2672_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1350_update_completed_
      -- 
    ca_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1350_inst_ack_1, ack => maxPool3D_CP_2672_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_sample_completed_
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1359_inst_ack_0, ack => maxPool3D_CP_2672_elements(6)); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(6), ack => RPIPE_maxpool_input_pipe_1359_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1359_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Sample/$entry
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1359_inst_ack_1, ack => maxPool3D_CP_2672_elements(7)); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(7), ack => type_cast_1363_inst_req_0); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(7), ack => RPIPE_maxpool_input_pipe_1371_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_sample_completed_
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_0, ack => maxPool3D_CP_2672_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1363_update_completed_
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_1, ack => maxPool3D_CP_2672_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Sample/$exit
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1371_inst_ack_0, ack => maxPool3D_CP_2672_elements(10)); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(10), ack => RPIPE_maxpool_input_pipe_1371_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1371_update_completed_
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1371_inst_ack_1, ack => maxPool3D_CP_2672_elements(11)); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(11), ack => type_cast_1375_inst_req_0); -- 
    rr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(11), ack => RPIPE_maxpool_input_pipe_1384_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Sample/$exit
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_0, ack => maxPool3D_CP_2672_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	50 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1375_update_completed_
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1375_inst_ack_1, ack => maxPool3D_CP_2672_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Sample/$exit
      -- 
    ra_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_0, ack => maxPool3D_CP_2672_elements(14)); -- 
    cr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(14), ack => RPIPE_maxpool_input_pipe_1384_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1384_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Sample/$entry
      -- 
    ca_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_1, ack => maxPool3D_CP_2672_elements(15)); -- 
    rr_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(15), ack => type_cast_1388_inst_req_0); -- 
    rr_2844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(15), ack => RPIPE_maxpool_input_pipe_1396_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Sample/$exit
      -- 
    ra_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => maxPool3D_CP_2672_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	50 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1388_update_completed_
      -- 
    ca_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => maxPool3D_CP_2672_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_update_start_
      -- 
    ra_2845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1396_inst_ack_0, ack => maxPool3D_CP_2672_elements(18)); -- 
    cr_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(18), ack => RPIPE_maxpool_input_pipe_1396_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1396_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Sample/rr
      -- 
    ca_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1396_inst_ack_1, ack => maxPool3D_CP_2672_elements(19)); -- 
    rr_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(19), ack => type_cast_1400_inst_req_0); -- 
    rr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(19), ack => RPIPE_maxpool_input_pipe_1409_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_sample_completed_
      -- 
    ra_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1400_inst_ack_0, ack => maxPool3D_CP_2672_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	50 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1400_Update/$exit
      -- 
    ca_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1400_inst_ack_1, ack => maxPool3D_CP_2672_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Update/cr
      -- 
    ra_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1409_inst_ack_0, ack => maxPool3D_CP_2672_elements(22)); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(22), ack => RPIPE_maxpool_input_pipe_1409_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1409_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Sample/rr
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1409_inst_ack_1, ack => maxPool3D_CP_2672_elements(23)); -- 
    rr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(23), ack => type_cast_1413_inst_req_0); -- 
    rr_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(23), ack => RPIPE_maxpool_input_pipe_1421_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Sample/ra
      -- 
    ra_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1413_inst_ack_0, ack => maxPool3D_CP_2672_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1413_Update/ca
      -- 
    ca_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1413_inst_ack_1, ack => maxPool3D_CP_2672_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Update/cr
      -- 
    ra_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1421_inst_ack_0, ack => maxPool3D_CP_2672_elements(26)); -- 
    cr_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(26), ack => RPIPE_maxpool_input_pipe_1421_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1421_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Sample/rr
      -- 
    ca_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1421_inst_ack_1, ack => maxPool3D_CP_2672_elements(27)); -- 
    rr_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(27), ack => type_cast_1425_inst_req_0); -- 
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(27), ack => RPIPE_maxpool_input_pipe_1434_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Sample/ra
      -- 
    ra_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => maxPool3D_CP_2672_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	50 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1425_Update/ca
      -- 
    ca_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => maxPool3D_CP_2672_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Update/cr
      -- 
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1434_inst_ack_0, ack => maxPool3D_CP_2672_elements(30)); -- 
    cr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(30), ack => RPIPE_maxpool_input_pipe_1434_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1434_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Sample/rr
      -- 
    ca_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1434_inst_ack_1, ack => maxPool3D_CP_2672_elements(31)); -- 
    rr_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(31), ack => type_cast_1438_inst_req_0); -- 
    rr_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(31), ack => RPIPE_maxpool_input_pipe_1446_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Sample/ra
      -- 
    ra_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_0, ack => maxPool3D_CP_2672_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	50 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1438_Update/ca
      -- 
    ca_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_1, ack => maxPool3D_CP_2672_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Update/cr
      -- 
    ra_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1446_inst_ack_0, ack => maxPool3D_CP_2672_elements(34)); -- 
    cr_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(34), ack => RPIPE_maxpool_input_pipe_1446_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1446_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Sample/rr
      -- 
    ca_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1446_inst_ack_1, ack => maxPool3D_CP_2672_elements(35)); -- 
    rr_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(35), ack => type_cast_1450_inst_req_0); -- 
    rr_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(35), ack => RPIPE_maxpool_input_pipe_1459_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Sample/ra
      -- 
    ra_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1450_inst_ack_0, ack => maxPool3D_CP_2672_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	50 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1450_Update/ca
      -- 
    ca_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1450_inst_ack_1, ack => maxPool3D_CP_2672_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Update/cr
      -- 
    ra_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1459_inst_ack_0, ack => maxPool3D_CP_2672_elements(38)); -- 
    cr_2989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(38), ack => RPIPE_maxpool_input_pipe_1459_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1459_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Sample/rr
      -- 
    ca_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1459_inst_ack_1, ack => maxPool3D_CP_2672_elements(39)); -- 
    rr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(39), ack => RPIPE_maxpool_input_pipe_1471_inst_req_0); -- 
    rr_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(39), ack => type_cast_1463_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Sample/ra
      -- 
    ra_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_0, ack => maxPool3D_CP_2672_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1463_Update/ca
      -- 
    ca_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1463_inst_ack_1, ack => maxPool3D_CP_2672_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Update/cr
      -- 
    ra_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1471_inst_ack_0, ack => maxPool3D_CP_2672_elements(42)); -- 
    cr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(42), ack => RPIPE_maxpool_input_pipe_1471_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1471_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Sample/rr
      -- 
    ca_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1471_inst_ack_1, ack => maxPool3D_CP_2672_elements(43)); -- 
    rr_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(43), ack => type_cast_1475_inst_req_0); -- 
    rr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(43), ack => RPIPE_maxpool_input_pipe_1484_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Sample/ra
      -- 
    ra_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1475_inst_ack_0, ack => maxPool3D_CP_2672_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1475_Update/ca
      -- 
    ca_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1475_inst_ack_1, ack => maxPool3D_CP_2672_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Update/cr
      -- 
    ra_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1484_inst_ack_0, ack => maxPool3D_CP_2672_elements(46)); -- 
    cr_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(46), ack => RPIPE_maxpool_input_pipe_1484_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/RPIPE_maxpool_input_pipe_1484_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Sample/rr
      -- 
    ca_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1484_inst_ack_1, ack => maxPool3D_CP_2672_elements(47)); -- 
    rr_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(47), ack => type_cast_1488_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Sample/ra
      -- 
    ra_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_0, ack => maxPool3D_CP_2672_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/type_cast_1488_Update/ca
      -- 
    ca_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_1, ack => maxPool3D_CP_2672_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	37 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	9 
    -- CP-element group 50: 	13 
    -- CP-element group 50: 	17 
    -- CP-element group 50: 	21 
    -- CP-element group 50: 	25 
    -- CP-element group 50: 	29 
    -- CP-element group 50: 	33 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515__entry__
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494__exit__
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1347_to_assign_stmt_1494/$exit
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/$entry
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Update/cr
      -- 
    rr_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(50), ack => type_cast_1498_inst_req_0); -- 
    cr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(50), ack => type_cast_1498_inst_req_1); -- 
    maxPool3D_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(37) & maxPool3D_CP_2672_elements(41) & maxPool3D_CP_2672_elements(45) & maxPool3D_CP_2672_elements(49) & maxPool3D_CP_2672_elements(5) & maxPool3D_CP_2672_elements(9) & maxPool3D_CP_2672_elements(13) & maxPool3D_CP_2672_elements(17) & maxPool3D_CP_2672_elements(21) & maxPool3D_CP_2672_elements(25) & maxPool3D_CP_2672_elements(29) & maxPool3D_CP_2672_elements(33);
      gj_maxPool3D_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Sample/ra
      -- 
    ra_3072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_0, ack => maxPool3D_CP_2672_elements(51)); -- 
    -- CP-element group 52:  branch  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (13) 
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516__entry__
      -- CP-element group 52: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515__exit__
      -- CP-element group 52: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/$exit
      -- CP-element group 52: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1344/assign_stmt_1499_to_assign_stmt_1515/type_cast_1498_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_dead_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_1344/R_cmp196_1517_place
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_if_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1344/if_stmt_1516_else_link/$entry
      -- 
    ca_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1498_inst_ack_1, ack => maxPool3D_CP_2672_elements(52)); -- 
    branch_req_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(52), ack => if_stmt_1516_branch_req_0); -- 
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (18) 
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567__entry__
      -- CP-element group 53: 	 branch_block_stmt_1344/merge_stmt_1522__exit__
      -- CP-element group 53: 	 branch_block_stmt_1344/if_stmt_1516_if_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1344/if_stmt_1516_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1344/entry_bbx_xnph
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/$entry
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1344/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1344/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1344/merge_stmt_1522_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_1344/merge_stmt_1522_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_1344/merge_stmt_1522_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_1344/merge_stmt_1522_PhiAck/dummy
      -- 
    if_choice_transition_3090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1516_branch_ack_1, ack => maxPool3D_CP_2672_elements(53)); -- 
    rr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(53), ack => type_cast_1553_inst_req_0); -- 
    cr_3112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(53), ack => type_cast_1553_inst_req_1); -- 
    -- CP-element group 54:  transition  place  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	204 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1344/if_stmt_1516_else_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_1344/if_stmt_1516_else_link/else_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_1344/entry_forx_xend
      -- CP-element group 54: 	 branch_block_stmt_1344/entry_forx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1344/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1516_branch_ack_0, ack => maxPool3D_CP_2672_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Sample/ra
      -- 
    ra_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_0, ack => maxPool3D_CP_2672_elements(55)); -- 
    -- CP-element group 56:  transition  place  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	198 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody
      -- CP-element group 56: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567__exit__
      -- CP-element group 56: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/$exit
      -- CP-element group 56: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1344/assign_stmt_1527_to_assign_stmt_1567/type_cast_1553_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/$entry
      -- CP-element group 56: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$entry
      -- 
    ca_3113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1553_inst_ack_1, ack => maxPool3D_CP_2672_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	203 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Sample/cra
      -- 
    cra_3125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1579_call_ack_0, ack => maxPool3D_CP_2672_elements(57)); -- 
    -- CP-element group 58:  branch  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	203 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591__entry__
      -- CP-element group 58: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590__exit__
      -- CP-element group 58: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/$exit
      -- CP-element group 58: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Update/cca
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1344/R_exitcond1_1592_place
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1344/if_stmt_1591_else_link/$entry
      -- 
    cca_3130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1579_call_ack_1, ack => maxPool3D_CP_2672_elements(58)); -- 
    branch_req_3138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(58), ack => if_stmt_1591_branch_req_0); -- 
    -- CP-element group 59:  merge  transition  place  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	204 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xendx_xloopexit_forx_xend
      -- CP-element group 59: 	 branch_block_stmt_1344/merge_stmt_1597__exit__
      -- CP-element group 59: 	 branch_block_stmt_1344/if_stmt_1591_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1344/if_stmt_1591_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1344/merge_stmt_1597_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1344/merge_stmt_1597_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1344/merge_stmt_1597_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1344/merge_stmt_1597_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1344/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1591_branch_ack_1, ack => maxPool3D_CP_2672_elements(59)); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	199 
    -- CP-element group 60: 	200 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_1344/if_stmt_1591_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1344/if_stmt_1591_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1591_branch_ack_0, ack => maxPool3D_CP_2672_elements(60)); -- 
    rr_3655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(60), ack => type_cast_1576_inst_req_0); -- 
    cr_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(60), ack => type_cast_1576_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	204 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Sample/cra
      -- 
    cra_3164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1614_call_ack_0, ack => maxPool3D_CP_2672_elements(61)); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	204 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	65 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	67 
    -- CP-element group 62: 	68 
    -- CP-element group 62:  members (25) 
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638__entry__
      -- CP-element group 62: 	 branch_block_stmt_1344/call_stmt_1614__exit__
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/call_stmt_1614/$exit
      -- CP-element group 62: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Update/cca
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Sample/rr
      -- 
    cca_3169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1614_call_ack_1, ack => maxPool3D_CP_2672_elements(62)); -- 
    cr_3199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1622_inst_req_1); -- 
    cr_3213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1626_inst_req_1); -- 
    rr_3208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1626_inst_req_0); -- 
    rr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1618_inst_req_0); -- 
    cr_3185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1618_inst_req_1); -- 
    rr_3194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(62), ack => type_cast_1622_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Sample/ra
      -- 
    ra_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_0, ack => maxPool3D_CP_2672_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1618_Update/ca
      -- 
    ca_3186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_1, ack => maxPool3D_CP_2672_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Sample/ra
      -- 
    ra_3195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1622_inst_ack_0, ack => maxPool3D_CP_2672_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1622_update_completed_
      -- 
    ca_3200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1622_inst_ack_1, ack => maxPool3D_CP_2672_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	62 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Sample/$exit
      -- 
    ra_3209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_0, ack => maxPool3D_CP_2672_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	62 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/type_cast_1626_update_completed_
      -- 
    ca_3214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_1, ack => maxPool3D_CP_2672_elements(68)); -- 
    -- CP-element group 69:  join  transition  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	66 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_1344/forx_xend_whilex_xbody
      -- CP-element group 69: 	 branch_block_stmt_1344/merge_stmt_1640__exit__
      -- CP-element group 69: 	 branch_block_stmt_1344/do_while_stmt_1657__entry__
      -- CP-element group 69: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638__exit__
      -- CP-element group 69: 	 branch_block_stmt_1344/assign_stmt_1619_to_assign_stmt_1638/$exit
      -- CP-element group 69: 	 branch_block_stmt_1344/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1344/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1344/merge_stmt_1640_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1344/merge_stmt_1640_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1344/merge_stmt_1640_PhiAck/$exit
      -- 
    maxPool3D_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(64) & maxPool3D_CP_2672_elements(66) & maxPool3D_CP_2672_elements(68);
      gj_maxPool3D_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  place  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	76 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1344/do_while_stmt_1657/$entry
      -- CP-element group 70: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657__entry__
      -- 
    maxPool3D_CP_2672_elements(70) <= maxPool3D_CP_2672_elements(69);
    -- CP-element group 71:  merge  place  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	180 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657__exit__
      -- 
    -- Element group maxPool3D_CP_2672_elements(71) is bound as output of CP function.
    -- CP-element group 72:  merge  place  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_back
      -- 
    -- Element group maxPool3D_CP_2672_elements(72) is bound as output of CP function.
    -- CP-element group 73:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	78 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	178 
    -- CP-element group 73: 	179 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_taken/$entry
      -- CP-element group 73: 	 branch_block_stmt_1344/do_while_stmt_1657/condition_done
      -- CP-element group 73: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_exit/$entry
      -- 
    maxPool3D_CP_2672_elements(73) <= maxPool3D_CP_2672_elements(78);
    -- CP-element group 74:  branch  place  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	177 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_body_done
      -- 
    maxPool3D_CP_2672_elements(74) <= maxPool3D_CP_2672_elements(177);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	87 
    -- CP-element group 75: 	108 
    -- CP-element group 75: 	129 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/back_edge_to_loop_body
      -- 
    maxPool3D_CP_2672_elements(75) <= maxPool3D_CP_2672_elements(72);
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	70 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	89 
    -- CP-element group 76: 	110 
    -- CP-element group 76: 	131 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/first_time_through_loop_body
      -- 
    maxPool3D_CP_2672_elements(76) <= maxPool3D_CP_2672_elements(70);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	103 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	176 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/loop_body_start
      -- CP-element group 77: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/$entry
      -- 
    -- Element group maxPool3D_CP_2672_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	171 
    -- CP-element group 78: 	175 
    -- CP-element group 78: 	176 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	73 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/condition_evaluated
      -- 
    condition_evaluated_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(78), ack => do_while_stmt_1657_branch_req_0); -- 
    maxPool3D_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(82) & maxPool3D_CP_2672_elements(171) & maxPool3D_CP_2672_elements(175) & maxPool3D_CP_2672_elements(176);
      gj_maxPool3D_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	102 
    -- CP-element group 79: 	123 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	104 
    -- CP-element group 79: 	125 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_sample_start__ps
      -- CP-element group 79: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/aggregated_phi_sample_req
      -- 
    maxPool3D_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(83) & maxPool3D_CP_2672_elements(102) & maxPool3D_CP_2672_elements(123) & maxPool3D_CP_2672_elements(82);
      gj_maxPool3D_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	85 
    -- CP-element group 80: 	105 
    -- CP-element group 80: 	126 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	161 
    -- CP-element group 80: 	165 
    -- CP-element group 80: 	169 
    -- CP-element group 80: 	173 
    -- CP-element group 80: 	177 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80: 	102 
    -- CP-element group 80: 	123 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/aggregated_phi_sample_ack
      -- 
    maxPool3D_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(85) & maxPool3D_CP_2672_elements(105) & maxPool3D_CP_2672_elements(126);
      gj_maxPool3D_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: 	103 
    -- CP-element group 81: 	124 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	106 
    -- CP-element group 81: 	127 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_update_start__ps
      -- CP-element group 81: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/aggregated_phi_update_req
      -- 
    maxPool3D_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(84) & maxPool3D_CP_2672_elements(103) & maxPool3D_CP_2672_elements(124);
      gj_maxPool3D_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	86 
    -- CP-element group 82: 	107 
    -- CP-element group 82: 	128 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/aggregated_phi_update_ack
      -- 
    maxPool3D_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(86) & maxPool3D_CP_2672_elements(107) & maxPool3D_CP_2672_elements(128);
      gj_maxPool3D_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	171 
    -- CP-element group 83: 	175 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_sample_start_
      -- 
    maxPool3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(171) & maxPool3D_CP_2672_elements(175);
      gj_maxPool3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: 	154 
    -- CP-element group 84: 	174 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	81 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_update_start_
      -- 
    maxPool3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(86) & maxPool3D_CP_2672_elements(154) & maxPool3D_CP_2672_elements(174);
      gj_maxPool3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	80 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	152 
    -- CP-element group 86: 	172 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(86) is bound as output of CP function.
    -- CP-element group 87:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	75 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_loopback_trigger
      -- 
    maxPool3D_CP_2672_elements(87) <= maxPool3D_CP_2672_elements(75);
    -- CP-element group 88:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_loopback_sample_req
      -- CP-element group 88: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_loopback_sample_req_ps
      -- 
    phi_stmt_1659_loopback_sample_req_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1659_loopback_sample_req_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(88), ack => phi_stmt_1659_req_0); -- 
    -- Element group maxPool3D_CP_2672_elements(88) is bound as output of CP function.
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	76 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_entry_trigger
      -- 
    maxPool3D_CP_2672_elements(89) <= maxPool3D_CP_2672_elements(76);
    -- CP-element group 90:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_entry_sample_req
      -- CP-element group 90: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_entry_sample_req_ps
      -- 
    phi_stmt_1659_entry_sample_req_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1659_entry_sample_req_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(90), ack => phi_stmt_1659_req_1); -- 
    -- Element group maxPool3D_CP_2672_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_phi_mux_ack_ps
      -- CP-element group 91: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1659_phi_mux_ack
      -- 
    phi_stmt_1659_phi_mux_ack_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1659_ack_0, ack => maxPool3D_CP_2672_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_sample_start_
      -- 
    rr_3263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(94), ack => type_cast_1662_inst_req_0); -- 
    maxPool3D_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(92) & maxPool3D_CP_2672_elements(96);
      gj_maxPool3D_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_update_start_
      -- 
    cr_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(95), ack => type_cast_1662_inst_req_1); -- 
    maxPool3D_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(93) & maxPool3D_CP_2672_elements(97);
      gj_maxPool3D_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_sample_completed_
      -- 
    ra_3264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_0, ack => maxPool3D_CP_2672_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1662_update_completed__ps
      -- 
    ca_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1662_inst_ack_1, ack => maxPool3D_CP_2672_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_update_completed__ps
      -- 
    maxPool3D_CP_2672_elements(100) <= maxPool3D_CP_2672_elements(101);
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	100 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_rowx_x1_at_entry_1663_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => maxPool3D_CP_2672_elements(99), ack => maxPool3D_CP_2672_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	80 
    -- CP-element group 102: 	163 
    -- CP-element group 102: 	167 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	79 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_sample_start_
      -- 
    maxPool3D_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(163) & maxPool3D_CP_2672_elements(167);
      gj_maxPool3D_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	77 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	107 
    -- CP-element group 103: 	150 
    -- CP-element group 103: 	166 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	81 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_update_start_
      -- 
    maxPool3D_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(107) & maxPool3D_CP_2672_elements(150) & maxPool3D_CP_2672_elements(166);
      gj_maxPool3D_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	79 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_sample_start__ps
      -- 
    maxPool3D_CP_2672_elements(104) <= maxPool3D_CP_2672_elements(79);
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	80 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	81 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_update_start__ps
      -- 
    maxPool3D_CP_2672_elements(106) <= maxPool3D_CP_2672_elements(81);
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	82 
    -- CP-element group 107: 	148 
    -- CP-element group 107: 	164 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	103 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	75 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_loopback_trigger
      -- 
    maxPool3D_CP_2672_elements(108) <= maxPool3D_CP_2672_elements(75);
    -- CP-element group 109:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_loopback_sample_req
      -- CP-element group 109: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_loopback_sample_req_ps
      -- 
    phi_stmt_1664_loopback_sample_req_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1664_loopback_sample_req_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(109), ack => phi_stmt_1664_req_0); -- 
    -- Element group maxPool3D_CP_2672_elements(109) is bound as output of CP function.
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_entry_trigger
      -- 
    maxPool3D_CP_2672_elements(110) <= maxPool3D_CP_2672_elements(76);
    -- CP-element group 111:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_entry_sample_req_ps
      -- CP-element group 111: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_entry_sample_req
      -- 
    phi_stmt_1664_entry_sample_req_3291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1664_entry_sample_req_3291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(111), ack => phi_stmt_1664_req_1); -- 
    -- Element group maxPool3D_CP_2672_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_phi_mux_ack_ps
      -- CP-element group 112: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1664_phi_mux_ack
      -- 
    phi_stmt_1664_phi_mux_ack_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1664_ack_0, ack => maxPool3D_CP_2672_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_sample_start_
      -- 
    rr_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(115), ack => type_cast_1667_inst_req_0); -- 
    maxPool3D_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(113) & maxPool3D_CP_2672_elements(117);
      gj_maxPool3D_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Update/$entry
      -- 
    cr_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(116), ack => type_cast_1667_inst_req_1); -- 
    maxPool3D_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(114) & maxPool3D_CP_2672_elements(118);
      gj_maxPool3D_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_sample_completed__ps
      -- 
    ra_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_0, ack => maxPool3D_CP_2672_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1667_Update/ca
      -- 
    ca_3313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1667_inst_ack_1, ack => maxPool3D_CP_2672_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_sample_completed__ps
      -- CP-element group 119: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_update_start_
      -- CP-element group 120: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_update_completed__ps
      -- 
    maxPool3D_CP_2672_elements(121) <= maxPool3D_CP_2672_elements(122);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	121 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_colx_x1_at_entry_1668_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => maxPool3D_CP_2672_elements(120), ack => maxPool3D_CP_2672_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	80 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	79 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_sample_start_
      -- 
    maxPool3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(80);
      gj_maxPool3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	146 
    -- CP-element group 124: 	162 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	81 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_update_start_
      -- 
    maxPool3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(77) & maxPool3D_CP_2672_elements(128) & maxPool3D_CP_2672_elements(146) & maxPool3D_CP_2672_elements(162);
      gj_maxPool3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_sample_start__ps
      -- 
    maxPool3D_CP_2672_elements(125) <= maxPool3D_CP_2672_elements(79);
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	80 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(126) is bound as output of CP function.
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	81 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_update_start__ps
      -- 
    maxPool3D_CP_2672_elements(127) <= maxPool3D_CP_2672_elements(81);
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	82 
    -- CP-element group 128: 	144 
    -- CP-element group 128: 	160 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	124 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(128) is bound as output of CP function.
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	75 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_loopback_trigger
      -- 
    maxPool3D_CP_2672_elements(129) <= maxPool3D_CP_2672_elements(75);
    -- CP-element group 130:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_loopback_sample_req_ps
      -- CP-element group 130: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_loopback_sample_req
      -- 
    phi_stmt_1669_loopback_sample_req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1669_loopback_sample_req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(130), ack => phi_stmt_1669_req_0); -- 
    -- Element group maxPool3D_CP_2672_elements(130) is bound as output of CP function.
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	76 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_entry_trigger
      -- 
    maxPool3D_CP_2672_elements(131) <= maxPool3D_CP_2672_elements(76);
    -- CP-element group 132:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_entry_sample_req_ps
      -- CP-element group 132: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_entry_sample_req
      -- 
    phi_stmt_1669_entry_sample_req_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1669_entry_sample_req_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(132), ack => phi_stmt_1669_req_1); -- 
    -- Element group maxPool3D_CP_2672_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_phi_mux_ack_ps
      -- CP-element group 133: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/phi_stmt_1669_phi_mux_ack
      -- 
    phi_stmt_1669_phi_mux_ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1669_ack_0, ack => maxPool3D_CP_2672_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2672_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_sample_start_
      -- 
    rr_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(136), ack => type_cast_1672_inst_req_0); -- 
    maxPool3D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(134) & maxPool3D_CP_2672_elements(138);
      gj_maxPool3D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_update_start_
      -- 
    cr_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(137), ack => type_cast_1672_inst_req_1); -- 
    maxPool3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(135) & maxPool3D_CP_2672_elements(139);
      gj_maxPool3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_sample_completed__ps
      -- 
    ra_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_0, ack => maxPool3D_CP_2672_elements(138)); -- 
    -- CP-element group 139:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1672_update_completed__ps
      -- 
    ca_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_1, ack => maxPool3D_CP_2672_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_sample_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_update_start_
      -- 
    -- Element group maxPool3D_CP_2672_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_update_completed__ps
      -- 
    maxPool3D_CP_2672_elements(142) <= maxPool3D_CP_2672_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/R_chlx_x0_at_entry_1673_update_completed_
      -- 
    -- Element group maxPool3D_CP_2672_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => maxPool3D_CP_2672_elements(141), ack => maxPool3D_CP_2672_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	128 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Sample/$entry
      -- 
    rr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(144), ack => type_cast_1677_inst_req_0); -- 
    maxPool3D_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(128) & maxPool3D_CP_2672_elements(146);
      gj_maxPool3D_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	158 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_update_start_
      -- 
    cr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(145), ack => type_cast_1677_inst_req_1); -- 
    maxPool3D_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(147) & maxPool3D_CP_2672_elements(158);
      gj_maxPool3D_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	124 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_sample_completed_
      -- 
    ra_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_0, ack => maxPool3D_CP_2672_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	156 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1677_update_completed_
      -- 
    ca_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1677_inst_ack_1, ack => maxPool3D_CP_2672_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	107 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_sample_start_
      -- 
    rr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(148), ack => type_cast_1681_inst_req_0); -- 
    maxPool3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(107) & maxPool3D_CP_2672_elements(150);
      gj_maxPool3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	158 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_update_start_
      -- 
    cr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(149), ack => type_cast_1681_inst_req_1); -- 
    maxPool3D_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(151) & maxPool3D_CP_2672_elements(158);
      gj_maxPool3D_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	103 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_sample_completed_
      -- 
    ra_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_0, ack => maxPool3D_CP_2672_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1681_update_completed_
      -- 
    ca_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1681_inst_ack_1, ack => maxPool3D_CP_2672_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	86 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Sample/rr
      -- 
    rr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(152), ack => type_cast_1685_inst_req_0); -- 
    maxPool3D_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(86) & maxPool3D_CP_2672_elements(154);
      gj_maxPool3D_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	158 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_update_start_
      -- CP-element group 153: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Update/$entry
      -- 
    cr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(153), ack => type_cast_1685_inst_req_1); -- 
    maxPool3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(155) & maxPool3D_CP_2672_elements(158);
      gj_maxPool3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	84 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Sample/$exit
      -- 
    ra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1685_inst_ack_0, ack => maxPool3D_CP_2672_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1685_Update/$exit
      -- 
    ca_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1685_inst_ack_1, ack => maxPool3D_CP_2672_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	147 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	155 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Sample/crr
      -- CP-element group 156: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_sample_start_
      -- 
    crr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(156), ack => call_stmt_1754_call_req_0); -- 
    maxPool3D_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(147) & maxPool3D_CP_2672_elements(151) & maxPool3D_CP_2672_elements(155) & maxPool3D_CP_2672_elements(158);
      gj_maxPool3D_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Update/ccr
      -- CP-element group 157: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_update_start_
      -- 
    ccr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(157), ack => call_stmt_1754_call_req_1); -- 
    maxPool3D_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_2672_elements(159);
      gj_maxPool3D_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: 	149 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Sample/cra
      -- CP-element group 158: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_sample_completed_
      -- 
    cra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1754_call_ack_0, ack => maxPool3D_CP_2672_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	177 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Update/cca
      -- CP-element group 159: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/call_stmt_1754_update_completed_
      -- 
    cca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1754_call_ack_1, ack => maxPool3D_CP_2672_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	128 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Sample/rr
      -- CP-element group 160: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_sample_start_
      -- 
    rr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(160), ack => type_cast_1768_inst_req_0); -- 
    maxPool3D_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(128) & maxPool3D_CP_2672_elements(162);
      gj_maxPool3D_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	80 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	170 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Update/cr
      -- CP-element group 161: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_update_start_
      -- CP-element group 161: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Update/$entry
      -- 
    cr_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(161), ack => type_cast_1768_inst_req_1); -- 
    maxPool3D_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(163) & maxPool3D_CP_2672_elements(170);
      gj_maxPool3D_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	124 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Sample/ra
      -- 
    ra_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_0, ack => maxPool3D_CP_2672_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	168 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	102 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1768_Update/$exit
      -- 
    ca_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_1, ack => maxPool3D_CP_2672_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	107 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Sample/req
      -- CP-element group 164: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_sample_start_
      -- 
    req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(164), ack => W_colx_x1_1760_delayed_1_0_1770_inst_req_0); -- 
    maxPool3D_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(107) & maxPool3D_CP_2672_elements(166);
      gj_maxPool3D_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	80 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	170 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_update_start_
      -- CP-element group 165: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Update/req
      -- CP-element group 165: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Update/$entry
      -- 
    req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(165), ack => W_colx_x1_1760_delayed_1_0_1770_inst_req_1); -- 
    maxPool3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(167) & maxPool3D_CP_2672_elements(170);
      gj_maxPool3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	103 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Sample/ack
      -- 
    ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1760_delayed_1_0_1770_inst_ack_0, ack => maxPool3D_CP_2672_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	102 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Update/ack
      -- CP-element group 167: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1772_Update/$exit
      -- 
    ack_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1760_delayed_1_0_1770_inst_ack_1, ack => maxPool3D_CP_2672_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	163 
    -- CP-element group 168: 	167 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_sample_start_
      -- 
    rr_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(168), ack => type_cast_1792_inst_req_0); -- 
    maxPool3D_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(163) & maxPool3D_CP_2672_elements(167) & maxPool3D_CP_2672_elements(170);
      gj_maxPool3D_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	80 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Update/cr
      -- CP-element group 169: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Update/$entry
      -- CP-element group 169: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_update_start_
      -- 
    cr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(169), ack => type_cast_1792_inst_req_1); -- 
    maxPool3D_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(171);
      gj_maxPool3D_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	161 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_sample_completed_
      -- 
    ra_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1792_inst_ack_0, ack => maxPool3D_CP_2672_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	78 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	83 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/type_cast_1792_update_completed_
      -- 
    ca_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1792_inst_ack_1, ack => maxPool3D_CP_2672_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	86 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Sample/req
      -- CP-element group 172: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_sample_start_
      -- 
    req_3472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(172), ack => W_rowx_x1_1781_delayed_2_0_1794_inst_req_0); -- 
    maxPool3D_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(86) & maxPool3D_CP_2672_elements(174);
      gj_maxPool3D_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	80 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Update/req
      -- CP-element group 173: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_update_start_
      -- 
    req_3477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(173), ack => W_rowx_x1_1781_delayed_2_0_1794_inst_req_1); -- 
    maxPool3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(175);
      gj_maxPool3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	84 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Sample/ack
      -- CP-element group 174: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_sample_completed_
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1781_delayed_2_0_1794_inst_ack_0, ack => maxPool3D_CP_2672_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	78 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	83 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/assign_stmt_1796_Update/ack
      -- 
    ack_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1781_delayed_2_0_1794_inst_ack_1, ack => maxPool3D_CP_2672_elements(175)); -- 
    -- CP-element group 176:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	77 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	78 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group maxPool3D_CP_2672_elements(176) is a control-delay.
    cp_element_176_delay: control_delay_element  generic map(name => " 176_delay", delay_value => 1)  port map(req => maxPool3D_CP_2672_elements(77), ack => maxPool3D_CP_2672_elements(176), clk => clk, reset =>reset);
    -- CP-element group 177:  join  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	80 
    -- CP-element group 177: 	159 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	74 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_1344/do_while_stmt_1657/do_while_stmt_1657_loop_body/$exit
      -- 
    maxPool3D_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(80) & maxPool3D_CP_2672_elements(159);
      gj_maxPool3D_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	73 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_exit/ack
      -- CP-element group 178: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_exit/$exit
      -- 
    ack_3483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1657_branch_ack_0, ack => maxPool3D_CP_2672_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	73 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_taken/ack
      -- CP-element group 179: 	 branch_block_stmt_1344/do_while_stmt_1657/loop_taken/$exit
      -- 
    ack_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1657_branch_ack_1, ack => maxPool3D_CP_2672_elements(179)); -- 
    -- CP-element group 180:  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	71 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	1 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_1344/do_while_stmt_1657/$exit
      -- 
    maxPool3D_CP_2672_elements(180) <= maxPool3D_CP_2672_elements(71);
    -- CP-element group 181:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	1 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	184 
    -- CP-element group 181:  members (18) 
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830__entry__
      -- CP-element group 181: 	 branch_block_stmt_1344/merge_stmt_1824__exit__
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/$entry
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_update_start_
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_1344/whilex_xbody_whilex_xend
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_1344/if_stmt_1820_if_link/if_choice_transition
      -- CP-element group 181: 	 branch_block_stmt_1344/if_stmt_1820_if_link/$exit
      -- CP-element group 181: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1344/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_1344/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 181: 	 branch_block_stmt_1344/merge_stmt_1824_PhiReqMerge
      -- CP-element group 181: 	 branch_block_stmt_1344/merge_stmt_1824_PhiAck/$entry
      -- CP-element group 181: 	 branch_block_stmt_1344/merge_stmt_1824_PhiAck/$exit
      -- CP-element group 181: 	 branch_block_stmt_1344/merge_stmt_1824_PhiAck/dummy
      -- 
    if_choice_transition_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1820_branch_ack_1, ack => maxPool3D_CP_2672_elements(181)); -- 
    cr_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(181), ack => type_cast_1829_inst_req_1); -- 
    rr_3517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(181), ack => type_cast_1829_inst_req_0); -- 
    -- CP-element group 182:  merge  transition  place  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	1 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_1344/merge_stmt_1824__entry__
      -- CP-element group 182: 	 branch_block_stmt_1344/if_stmt_1820__exit__
      -- CP-element group 182: 	 branch_block_stmt_1344/if_stmt_1820_else_link/else_choice_transition
      -- CP-element group 182: 	 branch_block_stmt_1344/if_stmt_1820_else_link/$exit
      -- CP-element group 182: 	 branch_block_stmt_1344/merge_stmt_1824_dead_link/$entry
      -- 
    else_choice_transition_3505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1820_branch_ack_0, ack => maxPool3D_CP_2672_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Sample/$exit
      -- 
    ra_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_0, ack => maxPool3D_CP_2672_elements(183)); -- 
    -- CP-element group 184:  fork  transition  place  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	181 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	186 
    -- CP-element group 184: 	188 
    -- CP-element group 184:  members (16) 
      -- CP-element group 184: 	 branch_block_stmt_1344/assign_stmt_1830__exit__
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846__entry__
      -- CP-element group 184: 	 branch_block_stmt_1344/assign_stmt_1830/$exit
      -- CP-element group 184: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Update/ccr
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/$entry
      -- CP-element group 184: 	 branch_block_stmt_1344/assign_stmt_1830/type_cast_1829_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Sample/crr
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Update/cr
      -- 
    ca_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_1, ack => maxPool3D_CP_2672_elements(184)); -- 
    ccr_3539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(184), ack => call_stmt_1833_call_req_1); -- 
    crr_3534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(184), ack => call_stmt_1833_call_req_0); -- 
    cr_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(184), ack => type_cast_1837_inst_req_1); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Sample/cra
      -- CP-element group 185: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Sample/$exit
      -- 
    cra_3535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1833_call_ack_0, ack => maxPool3D_CP_2672_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Update/cca
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/call_stmt_1833_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Sample/$entry
      -- 
    cca_3540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1833_call_ack_1, ack => maxPool3D_CP_2672_elements(186)); -- 
    rr_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(186), ack => type_cast_1837_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Sample/$exit
      -- 
    ra_3549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_0, ack => maxPool3D_CP_2672_elements(187)); -- 
    -- CP-element group 188:  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	184 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (6) 
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/type_cast_1837_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Sample/req
      -- 
    ca_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_1, ack => maxPool3D_CP_2672_elements(188)); -- 
    req_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(188), ack => WPIPE_elapsed_time_pipe_1844_inst_req_0); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_update_start_
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Sample/ack
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Update/req
      -- 
    ack_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1844_inst_ack_0, ack => maxPool3D_CP_2672_elements(189)); -- 
    req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(189), ack => WPIPE_elapsed_time_pipe_1844_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  place  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	193 
    -- CP-element group 190: 	194 
    -- CP-element group 190: 	197 
    -- CP-element group 190:  members (22) 
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867__entry__
      -- CP-element group 190: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846__exit__
      -- CP-element group 190: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/$exit
      -- CP-element group 190: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1344/call_stmt_1833_to_assign_stmt_1846/WPIPE_elapsed_time_pipe_1844_Update/ack
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_update_start_
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_update_start_
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_update_start_
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Update/ccr
      -- 
    ack_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1844_inst_ack_1, ack => maxPool3D_CP_2672_elements(190)); -- 
    rr_3579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(190), ack => type_cast_1850_inst_req_0); -- 
    cr_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(190), ack => type_cast_1850_inst_req_1); -- 
    rr_3593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(190), ack => type_cast_1854_inst_req_0); -- 
    cr_3598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(190), ack => type_cast_1854_inst_req_1); -- 
    ccr_3612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(190), ack => call_stmt_1867_call_req_1); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Sample/ra
      -- 
    ra_3580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_0, ack => maxPool3D_CP_2672_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1850_Update/ca
      -- 
    ca_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_1, ack => maxPool3D_CP_2672_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Sample/ra
      -- 
    ra_3594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1854_inst_ack_0, ack => maxPool3D_CP_2672_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/type_cast_1854_Update/ca
      -- 
    ca_3599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1854_inst_ack_1, ack => maxPool3D_CP_2672_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Sample/crr
      -- 
    crr_3607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(195), ack => call_stmt_1867_call_req_0); -- 
    maxPool3D_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(192) & maxPool3D_CP_2672_elements(194);
      gj_maxPool3D_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Sample/cra
      -- 
    cra_3608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1867_call_ack_0, ack => maxPool3D_CP_2672_elements(196)); -- 
    -- CP-element group 197:  transition  place  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	190 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (16) 
      -- CP-element group 197: 	 branch_block_stmt_1344/$exit
      -- CP-element group 197: 	 $exit
      -- CP-element group 197: 	 branch_block_stmt_1344/branch_block_stmt_1344__exit__
      -- CP-element group 197: 	 branch_block_stmt_1344/merge_stmt_1869__exit__
      -- CP-element group 197: 	 branch_block_stmt_1344/return__
      -- CP-element group 197: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867__exit__
      -- CP-element group 197: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/$exit
      -- CP-element group 197: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_1344/assign_stmt_1851_to_call_stmt_1867/call_stmt_1867_Update/cca
      -- CP-element group 197: 	 branch_block_stmt_1344/return___PhiReq/$entry
      -- CP-element group 197: 	 branch_block_stmt_1344/return___PhiReq/$exit
      -- CP-element group 197: 	 branch_block_stmt_1344/merge_stmt_1869_PhiReqMerge
      -- CP-element group 197: 	 branch_block_stmt_1344/merge_stmt_1869_PhiAck/$entry
      -- CP-element group 197: 	 branch_block_stmt_1344/merge_stmt_1869_PhiAck/$exit
      -- CP-element group 197: 	 branch_block_stmt_1344/merge_stmt_1869_PhiAck/dummy
      -- 
    cca_3613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1867_call_ack_1, ack => maxPool3D_CP_2672_elements(197)); -- 
    -- CP-element group 198:  transition  output  delay-element  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	56 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	202 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 198: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/$exit
      -- CP-element group 198: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$exit
      -- CP-element group 198: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1574_konst_delay_trans
      -- CP-element group 198: 	 branch_block_stmt_1344/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_req
      -- 
    phi_stmt_1570_req_3636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1570_req_3636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(198), ack => phi_stmt_1570_req_0); -- 
    -- Element group maxPool3D_CP_2672_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => maxPool3D_CP_2672_elements(56), ack => maxPool3D_CP_2672_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	60 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Sample/ra
      -- 
    ra_3656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1576_inst_ack_0, ack => maxPool3D_CP_2672_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	60 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (2) 
      -- CP-element group 200: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/Update/ca
      -- 
    ca_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1576_inst_ack_1, ack => maxPool3D_CP_2672_elements(200)); -- 
    -- CP-element group 201:  join  transition  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/$exit
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$exit
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/$exit
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1576/SplitProtocol/$exit
      -- CP-element group 201: 	 branch_block_stmt_1344/forx_xbody_forx_xbody_PhiReq/phi_stmt_1570/phi_stmt_1570_req
      -- 
    phi_stmt_1570_req_3662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1570_req_3662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(201), ack => phi_stmt_1570_req_1); -- 
    maxPool3D_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2672_elements(199) & maxPool3D_CP_2672_elements(200);
      gj_maxPool3D_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2672_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  merge  transition  place  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	198 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_1344/merge_stmt_1569_PhiReqMerge
      -- CP-element group 202: 	 branch_block_stmt_1344/merge_stmt_1569_PhiAck/$entry
      -- 
    maxPool3D_CP_2672_elements(202) <= OrReduce(maxPool3D_CP_2672_elements(198) & maxPool3D_CP_2672_elements(201));
    -- CP-element group 203:  fork  transition  place  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	57 
    -- CP-element group 203: 	58 
    -- CP-element group 203:  members (11) 
      -- CP-element group 203: 	 branch_block_stmt_1344/merge_stmt_1569__exit__
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590__entry__
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/$entry
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_update_start_
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Sample/crr
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_1344/call_stmt_1579_to_assign_stmt_1590/call_stmt_1579_Update/ccr
      -- CP-element group 203: 	 branch_block_stmt_1344/merge_stmt_1569_PhiAck/$exit
      -- CP-element group 203: 	 branch_block_stmt_1344/merge_stmt_1569_PhiAck/phi_stmt_1570_ack
      -- 
    phi_stmt_1570_ack_3667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1570_ack_0, ack => maxPool3D_CP_2672_elements(203)); -- 
    crr_3124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(203), ack => call_stmt_1579_call_req_0); -- 
    ccr_3129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(203), ack => call_stmt_1579_call_req_1); -- 
    -- CP-element group 204:  merge  fork  transition  place  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	54 
    -- CP-element group 204: 	59 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	61 
    -- CP-element group 204: 	62 
    -- CP-element group 204:  members (17) 
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614__entry__
      -- CP-element group 204: 	 branch_block_stmt_1344/assign_stmt_1606_to_assign_stmt_1611__exit__
      -- CP-element group 204: 	 branch_block_stmt_1344/assign_stmt_1606_to_assign_stmt_1611__entry__
      -- CP-element group 204: 	 branch_block_stmt_1344/merge_stmt_1599__exit__
      -- CP-element group 204: 	 branch_block_stmt_1344/assign_stmt_1606_to_assign_stmt_1611/$entry
      -- CP-element group 204: 	 branch_block_stmt_1344/assign_stmt_1606_to_assign_stmt_1611/$exit
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/$entry
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_update_start_
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Sample/crr
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_1344/call_stmt_1614/call_stmt_1614_Update/ccr
      -- CP-element group 204: 	 branch_block_stmt_1344/merge_stmt_1599_PhiReqMerge
      -- CP-element group 204: 	 branch_block_stmt_1344/merge_stmt_1599_PhiAck/$entry
      -- CP-element group 204: 	 branch_block_stmt_1344/merge_stmt_1599_PhiAck/$exit
      -- CP-element group 204: 	 branch_block_stmt_1344/merge_stmt_1599_PhiAck/dummy
      -- 
    crr_3163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(204), ack => call_stmt_1614_call_req_0); -- 
    ccr_3168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2672_elements(204), ack => call_stmt_1614_call_req_1); -- 
    maxPool3D_CP_2672_elements(204) <= OrReduce(maxPool3D_CP_2672_elements(54) & maxPool3D_CP_2672_elements(59));
    maxPool3D_do_while_stmt_1657_terminator_3488: loop_terminator -- 
      generic map (name => " maxPool3D_do_while_stmt_1657_terminator_3488", max_iterations_in_flight =>15) 
      port map(loop_body_exit => maxPool3D_CP_2672_elements(74),loop_continue => maxPool3D_CP_2672_elements(179),loop_terminate => maxPool3D_CP_2672_elements(178),loop_back => maxPool3D_CP_2672_elements(72),loop_exit => maxPool3D_CP_2672_elements(71),clk => clk, reset => reset); -- 
    phi_stmt_1659_phi_seq_3278_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2672_elements(87);
      maxPool3D_CP_2672_elements(92)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2672_elements(96);
      maxPool3D_CP_2672_elements(93)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2672_elements(97);
      maxPool3D_CP_2672_elements(88) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2672_elements(89);
      maxPool3D_CP_2672_elements(98)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2672_elements(98);
      maxPool3D_CP_2672_elements(99)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2672_elements(100);
      maxPool3D_CP_2672_elements(90) <= phi_mux_reqs(1);
      phi_stmt_1659_phi_seq_3278 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1659_phi_seq_3278") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2672_elements(79), 
          phi_sample_ack => maxPool3D_CP_2672_elements(85), 
          phi_update_req => maxPool3D_CP_2672_elements(81), 
          phi_update_ack => maxPool3D_CP_2672_elements(86), 
          phi_mux_ack => maxPool3D_CP_2672_elements(91), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1664_phi_seq_3322_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2672_elements(108);
      maxPool3D_CP_2672_elements(113)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2672_elements(117);
      maxPool3D_CP_2672_elements(114)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2672_elements(118);
      maxPool3D_CP_2672_elements(109) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2672_elements(110);
      maxPool3D_CP_2672_elements(119)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2672_elements(119);
      maxPool3D_CP_2672_elements(120)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2672_elements(121);
      maxPool3D_CP_2672_elements(111) <= phi_mux_reqs(1);
      phi_stmt_1664_phi_seq_3322 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1664_phi_seq_3322") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2672_elements(104), 
          phi_sample_ack => maxPool3D_CP_2672_elements(105), 
          phi_update_req => maxPool3D_CP_2672_elements(106), 
          phi_update_ack => maxPool3D_CP_2672_elements(107), 
          phi_mux_ack => maxPool3D_CP_2672_elements(112), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1669_phi_seq_3366_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2672_elements(129);
      maxPool3D_CP_2672_elements(134)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2672_elements(138);
      maxPool3D_CP_2672_elements(135)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2672_elements(139);
      maxPool3D_CP_2672_elements(130) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2672_elements(131);
      maxPool3D_CP_2672_elements(140)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2672_elements(140);
      maxPool3D_CP_2672_elements(141)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2672_elements(142);
      maxPool3D_CP_2672_elements(132) <= phi_mux_reqs(1);
      phi_stmt_1669_phi_seq_3366 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1669_phi_seq_3366") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2672_elements(125), 
          phi_sample_ack => maxPool3D_CP_2672_elements(126), 
          phi_update_req => maxPool3D_CP_2672_elements(127), 
          phi_update_ack => maxPool3D_CP_2672_elements(128), 
          phi_mux_ack => maxPool3D_CP_2672_elements(133), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3230_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= maxPool3D_CP_2672_elements(75);
        preds(1)  <= maxPool3D_CP_2672_elements(76);
        entry_tmerge_3230 : transition_merge -- 
          generic map(name => " entry_tmerge_3230")
          port map (preds => preds, symbol_out => maxPool3D_CP_2672_elements(77));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1819_wire : std_logic_vector(0 downto 0);
    signal add101_1638 : std_logic_vector(31 downto 0);
    signal add117_1696 : std_logic_vector(31 downto 0);
    signal add119_1706 : std_logic_vector(31 downto 0);
    signal add132_1722 : std_logic_vector(31 downto 0);
    signal add135_1732 : std_logic_vector(31 downto 0);
    signal add13_1394 : std_logic_vector(15 downto 0);
    signal add142_1737 : std_logic_vector(31 downto 0);
    signal add146_1742 : std_logic_vector(31 downto 0);
    signal add149_1747 : std_logic_vector(31 downto 0);
    signal add23_1419 : std_logic_vector(15 downto 0);
    signal add33_1444 : std_logic_vector(15 downto 0);
    signal add43_1469 : std_logic_vector(31 downto 0);
    signal add53_1494 : std_logic_vector(15 downto 0);
    signal add_1369 : std_logic_vector(31 downto 0);
    signal call11_1385 : std_logic_vector(7 downto 0);
    signal call150_1754 : std_logic_vector(7 downto 0);
    signal call16_1397 : std_logic_vector(7 downto 0);
    signal call180_1833 : std_logic_vector(63 downto 0);
    signal call21_1410 : std_logic_vector(7 downto 0);
    signal call26_1422 : std_logic_vector(7 downto 0);
    signal call2_1360 : std_logic_vector(7 downto 0);
    signal call31_1435 : std_logic_vector(7 downto 0);
    signal call36_1447 : std_logic_vector(7 downto 0);
    signal call41_1460 : std_logic_vector(7 downto 0);
    signal call46_1472 : std_logic_vector(7 downto 0);
    signal call51_1485 : std_logic_vector(7 downto 0);
    signal call6_1372 : std_logic_vector(7 downto 0);
    signal call89_1614 : std_logic_vector(63 downto 0);
    signal call_1347 : std_logic_vector(7 downto 0);
    signal chlx_x0_1669 : std_logic_vector(15 downto 0);
    signal chlx_x0_at_entry_1651 : std_logic_vector(15 downto 0);
    signal chlx_x1_1784 : std_logic_vector(15 downto 0);
    signal cmp157_1765 : std_logic_vector(0 downto 0);
    signal cmp165_1789 : std_logic_vector(0 downto 0);
    signal cmp175_1813 : std_logic_vector(0 downto 0);
    signal cmp196_1515 : std_logic_vector(0 downto 0);
    signal colx_x1_1664 : std_logic_vector(15 downto 0);
    signal colx_x1_1760_delayed_1_0_1772 : std_logic_vector(15 downto 0);
    signal colx_x1_at_entry_1646 : std_logic_vector(15 downto 0);
    signal colx_x2_1808 : std_logic_vector(15 downto 0);
    signal conv100_1623 : std_logic_vector(31 downto 0);
    signal conv107_1678 : std_logic_vector(31 downto 0);
    signal conv111_1682 : std_logic_vector(31 downto 0);
    signal conv113_1627 : std_logic_vector(31 downto 0);
    signal conv115_1686 : std_logic_vector(31 downto 0);
    signal conv12_1389 : std_logic_vector(15 downto 0);
    signal conv181_1838 : std_logic_vector(63 downto 0);
    signal conv189_1851 : std_logic_vector(31 downto 0);
    signal conv192_1855 : std_logic_vector(31 downto 0);
    signal conv19_1401 : std_logic_vector(15 downto 0);
    signal conv1_1351 : std_logic_vector(31 downto 0);
    signal conv22_1414 : std_logic_vector(15 downto 0);
    signal conv29_1426 : std_logic_vector(15 downto 0);
    signal conv32_1439 : std_logic_vector(15 downto 0);
    signal conv39_1451 : std_logic_vector(31 downto 0);
    signal conv3_1364 : std_logic_vector(31 downto 0);
    signal conv42_1464 : std_logic_vector(31 downto 0);
    signal conv49_1476 : std_logic_vector(15 downto 0);
    signal conv52_1489 : std_logic_vector(15 downto 0);
    signal conv59_1499 : std_logic_vector(31 downto 0);
    signal conv90_1830 : std_logic_vector(63 downto 0);
    signal conv98_1619 : std_logic_vector(31 downto 0);
    signal conv9_1376 : std_logic_vector(15 downto 0);
    signal exitcond1_1590 : std_logic_vector(0 downto 0);
    signal iNsTr_14_1554 : std_logic_vector(63 downto 0);
    signal iNsTr_20_1570 : std_logic_vector(63 downto 0);
    signal inc152_1760 : std_logic_vector(15 downto 0);
    signal inc160_1769 : std_logic_vector(15 downto 0);
    signal inc160x_xcolx_x1_1777 : std_logic_vector(15 downto 0);
    signal inc169_1793 : std_logic_vector(15 downto 0);
    signal inc169x_xrowx_x1_1801 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1585 : std_logic_vector(63 downto 0);
    signal mul116_1691 : std_logic_vector(31 downto 0);
    signal mul118_1701 : std_logic_vector(31 downto 0);
    signal mul131_1717 : std_logic_vector(31 downto 0);
    signal mul133_1633 : std_logic_vector(31 downto 0);
    signal mul190_1860 : std_logic_vector(31 downto 0);
    signal mul193_1865 : std_logic_vector(31 downto 0);
    signal mul62_1509 : std_logic_vector(31 downto 0);
    signal mul86_1611 : std_logic_vector(15 downto 0);
    signal mul_1504 : std_logic_vector(31 downto 0);
    signal rowx_x1_1659 : std_logic_vector(15 downto 0);
    signal rowx_x1_1781_delayed_2_0_1796 : std_logic_vector(15 downto 0);
    signal rowx_x1_at_entry_1641 : std_logic_vector(15 downto 0);
    signal shl10_1382 : std_logic_vector(15 downto 0);
    signal shl120_1712 : std_logic_vector(31 downto 0);
    signal shl134_1727 : std_logic_vector(31 downto 0);
    signal shl20_1407 : std_logic_vector(15 downto 0);
    signal shl30_1432 : std_logic_vector(15 downto 0);
    signal shl40_1457 : std_logic_vector(31 downto 0);
    signal shl50_1482 : std_logic_vector(15 downto 0);
    signal shl_1357 : std_logic_vector(31 downto 0);
    signal shr79194_1606 : std_logic_vector(15 downto 0);
    signal sub_1843 : std_logic_vector(63 downto 0);
    signal tmp199_1532 : std_logic_vector(31 downto 0);
    signal tmp200_1538 : std_logic_vector(31 downto 0);
    signal tmp200x_xop_1550 : std_logic_vector(31 downto 0);
    signal tmp201_1544 : std_logic_vector(0 downto 0);
    signal tmp204_1567 : std_logic_vector(63 downto 0);
    signal tmp_1527 : std_logic_vector(31 downto 0);
    signal type_cast_1355_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1405_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1455_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1480_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1542_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1548_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1565_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1574_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1576_wire : std_logic_vector(63 downto 0);
    signal type_cast_1583_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1631_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1662_wire : std_logic_vector(15 downto 0);
    signal type_cast_1667_wire : std_logic_vector(15 downto 0);
    signal type_cast_1672_wire : std_logic_vector(15 downto 0);
    signal type_cast_1710_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1758_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1781_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1805_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1828_wire : std_logic_vector(63 downto 0);
    signal type_cast_1836_wire : std_logic_vector(63 downto 0);
    signal whilex_xbody_whilex_xend_taken_1816 : std_logic_vector(0 downto 0);
    signal xx_xop_1560 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    chlx_x0_at_entry_1651 <= "0000000000000000";
    colx_x1_at_entry_1646 <= "0000000000000000";
    rowx_x1_at_entry_1641 <= "0000000000000000";
    type_cast_1355_wire_constant <= "00000000000000000000000000001000";
    type_cast_1380_wire_constant <= "0000000000001000";
    type_cast_1405_wire_constant <= "0000000000001000";
    type_cast_1430_wire_constant <= "0000000000001000";
    type_cast_1455_wire_constant <= "00000000000000000000000000001000";
    type_cast_1480_wire_constant <= "0000000000001000";
    type_cast_1513_wire_constant <= "00000000000000000000000000001111";
    type_cast_1536_wire_constant <= "00000000000000000000000000000100";
    type_cast_1542_wire_constant <= "00000000000000000000000000000001";
    type_cast_1548_wire_constant <= "11111111111111111111111111111111";
    type_cast_1558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1565_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1574_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1583_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1604_wire_constant <= "0000000000000100";
    type_cast_1631_wire_constant <= "00000000000000000000000000000001";
    type_cast_1710_wire_constant <= "00000000000000000000000000000010";
    type_cast_1758_wire_constant <= "0000000000000001";
    type_cast_1781_wire_constant <= "0000000000000000";
    type_cast_1805_wire_constant <= "0000000000000000";
    phi_stmt_1570: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1574_wire_constant & type_cast_1576_wire;
      req <= phi_stmt_1570_req_0 & phi_stmt_1570_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1570",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1570_ack_0,
          idata => idata,
          odata => iNsTr_20_1570,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1570
    phi_stmt_1659: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1662_wire & rowx_x1_at_entry_1641;
      req <= phi_stmt_1659_req_0 & phi_stmt_1659_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1659",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1659_ack_0,
          idata => idata,
          odata => rowx_x1_1659,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1659
    phi_stmt_1664: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1667_wire & colx_x1_at_entry_1646;
      req <= phi_stmt_1664_req_0 & phi_stmt_1664_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1664",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1664_ack_0,
          idata => idata,
          odata => colx_x1_1664,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1664
    phi_stmt_1669: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1672_wire & chlx_x0_at_entry_1651;
      req <= phi_stmt_1669_req_0 & phi_stmt_1669_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1669",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1669_ack_0,
          idata => idata,
          odata => chlx_x0_1669,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1669
    -- flow-through select operator MUX_1566_inst
    tmp204_1567 <= xx_xop_1560 when (tmp201_1544(0) /=  '0') else type_cast_1565_wire_constant;
    -- flow-through select operator MUX_1783_inst
    chlx_x1_1784 <= type_cast_1781_wire_constant when (cmp157_1765(0) /=  '0') else inc152_1760;
    -- flow-through select operator MUX_1807_inst
    colx_x2_1808 <= type_cast_1805_wire_constant when (cmp165_1789(0) /=  '0') else inc160x_xcolx_x1_1777;
    W_colx_x1_1760_delayed_1_0_1770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1_1760_delayed_1_0_1770_inst_req_0;
      W_colx_x1_1760_delayed_1_0_1770_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1_1760_delayed_1_0_1770_inst_req_1;
      W_colx_x1_1760_delayed_1_0_1770_inst_ack_1<= rack(0);
      W_colx_x1_1760_delayed_1_0_1770_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1_1760_delayed_1_0_1770_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1_1760_delayed_1_0_1772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rowx_x1_1781_delayed_2_0_1794_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rowx_x1_1781_delayed_2_0_1794_inst_req_0;
      W_rowx_x1_1781_delayed_2_0_1794_inst_ack_0<= wack(0);
      rreq(0) <= W_rowx_x1_1781_delayed_2_0_1794_inst_req_1;
      W_rowx_x1_1781_delayed_2_0_1794_inst_ack_1<= rack(0);
      W_rowx_x1_1781_delayed_2_0_1794_inst : InterlockBuffer generic map ( -- 
        name => "W_rowx_x1_1781_delayed_2_0_1794_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowx_x1_1781_delayed_2_0_1796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_1814_inst
    process(cmp175_1813) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp175_1813(0 downto 0);
      whilex_xbody_whilex_xend_taken_1816 <= tmp_var; -- 
    end process;
    type_cast_1350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1350_inst_req_0;
      type_cast_1350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1350_inst_req_1;
      type_cast_1350_inst_ack_1<= rack(0);
      type_cast_1350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1363_inst_req_0;
      type_cast_1363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1363_inst_req_1;
      type_cast_1363_inst_ack_1<= rack(0);
      type_cast_1363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1375_inst_req_0;
      type_cast_1375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1375_inst_req_1;
      type_cast_1375_inst_ack_1<= rack(0);
      type_cast_1375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1400_inst_req_0;
      type_cast_1400_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1400_inst_req_1;
      type_cast_1400_inst_ack_1<= rack(0);
      type_cast_1400_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1400_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1397,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1401,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1413_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1413_inst_req_0;
      type_cast_1413_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1413_inst_req_1;
      type_cast_1413_inst_ack_1<= rack(0);
      type_cast_1413_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1413_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1438_inst_req_0;
      type_cast_1438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1438_inst_req_1;
      type_cast_1438_inst_ack_1<= rack(0);
      type_cast_1438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1450_inst_req_0;
      type_cast_1450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1450_inst_req_1;
      type_cast_1450_inst_ack_1<= rack(0);
      type_cast_1450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1451,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1463_inst_req_0;
      type_cast_1463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1463_inst_req_1;
      type_cast_1463_inst_ack_1<= rack(0);
      type_cast_1463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1475_inst_req_0;
      type_cast_1475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1475_inst_req_1;
      type_cast_1475_inst_ack_1<= rack(0);
      type_cast_1475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1472,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1488_inst_req_0;
      type_cast_1488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1488_inst_req_1;
      type_cast_1488_inst_ack_1<= rack(0);
      type_cast_1488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1498_inst_req_0;
      type_cast_1498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1498_inst_req_1;
      type_cast_1498_inst_ack_1<= rack(0);
      type_cast_1498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1553_inst_req_0;
      type_cast_1553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1553_inst_req_1;
      type_cast_1553_inst_ack_1<= rack(0);
      type_cast_1553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp200x_xop_1550,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_1554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1576_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1576_inst_req_0;
      type_cast_1576_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1576_inst_req_1;
      type_cast_1576_inst_ack_1<= rack(0);
      type_cast_1576_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1576_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1576_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1618_inst_req_0;
      type_cast_1618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1618_inst_req_1;
      type_cast_1618_inst_ack_1<= rack(0);
      type_cast_1618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr79194_1606,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_1619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1622_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1622_inst_req_0;
      type_cast_1622_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1622_inst_req_1;
      type_cast_1622_inst_ack_1<= rack(0);
      type_cast_1622_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1622_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul86_1611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_1623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1626_inst_req_0;
      type_cast_1626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1626_inst_req_1;
      type_cast_1626_inst_ack_1<= rack(0);
      type_cast_1626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_1627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1662_inst_req_0;
      type_cast_1662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1662_inst_req_1;
      type_cast_1662_inst_ack_1<= rack(0);
      type_cast_1662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1662_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc169x_xrowx_x1_1801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1662_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1667_inst_req_0;
      type_cast_1667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1667_inst_req_1;
      type_cast_1667_inst_ack_1<= rack(0);
      type_cast_1667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1667_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2_1808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1667_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1672_inst_req_0;
      type_cast_1672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1672_inst_req_1;
      type_cast_1672_inst_ack_1<= rack(0);
      type_cast_1672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1672_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1_1784,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1672_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1677_inst_req_0;
      type_cast_1677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1677_inst_req_1;
      type_cast_1677_inst_ack_1<= rack(0);
      type_cast_1677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0_1669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1678,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1681_inst_req_0;
      type_cast_1681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1681_inst_req_1;
      type_cast_1681_inst_ack_1<= rack(0);
      type_cast_1681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1685_inst_req_0;
      type_cast_1685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1685_inst_req_1;
      type_cast_1685_inst_ack_1<= rack(0);
      type_cast_1685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1768_inst_req_0;
      type_cast_1768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1768_inst_req_1;
      type_cast_1768_inst_ack_1<= rack(0);
      type_cast_1768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1768_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp157_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc160_1769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1792_inst_req_0;
      type_cast_1792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1792_inst_req_1;
      type_cast_1792_inst_ack_1<= rack(0);
      type_cast_1792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1792_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp165_1789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc169_1793,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1829_inst_req_0;
      type_cast_1829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1829_inst_req_1;
      type_cast_1829_inst_ack_1<= rack(0);
      type_cast_1829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1828_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1837_inst_req_0;
      type_cast_1837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1837_inst_req_1;
      type_cast_1837_inst_ack_1<= rack(0);
      type_cast_1837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1836_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_1838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1850_inst_req_0;
      type_cast_1850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1850_inst_req_1;
      type_cast_1850_inst_ack_1<= rack(0);
      type_cast_1850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv189_1851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1854_inst_req_0;
      type_cast_1854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1854_inst_req_1;
      type_cast_1854_inst_ack_1<= rack(0);
      type_cast_1854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_1855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1657_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1819_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1657_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1657_branch_req_0,
          ack0 => do_while_stmt_1657_branch_ack_0,
          ack1 => do_while_stmt_1657_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1516_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp196_1515;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1516_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1516_branch_req_0,
          ack0 => if_stmt_1516_branch_ack_0,
          ack1 => if_stmt_1516_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1591_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1590;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1591_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1591_branch_req_0,
          ack0 => if_stmt_1591_branch_ack_0,
          ack1 => if_stmt_1591_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1820_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_1816;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1820_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1820_branch_req_0,
          ack0 => if_stmt_1820_branch_ack_0,
          ack1 => if_stmt_1820_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1759_inst
    process(chlx_x0_1669) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0_1669, type_cast_1758_wire_constant, tmp_var);
      inc152_1760 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1776_inst
    process(inc160_1769, colx_x1_1760_delayed_1_0_1772) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc160_1769, colx_x1_1760_delayed_1_0_1772, tmp_var);
      inc160x_xcolx_x1_1777 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1800_inst
    process(inc169_1793, rowx_x1_1781_delayed_2_0_1796) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc169_1793, rowx_x1_1781_delayed_2_0_1796, tmp_var);
      inc169x_xrowx_x1_1801 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1549_inst
    process(tmp200_1538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp200_1538, type_cast_1548_wire_constant, tmp_var);
      tmp200x_xop_1550 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1637_inst
    process(conv100_1623, conv98_1619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_1623, conv98_1619, tmp_var);
      add101_1638 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1695_inst
    process(conv111_1682, mul116_1691) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_1682, mul116_1691, tmp_var);
      add117_1696 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1705_inst
    process(mul118_1701, conv107_1678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul118_1701, conv107_1678, tmp_var);
      add119_1706 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1721_inst
    process(conv111_1682, mul131_1717) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_1682, mul131_1717, tmp_var);
      add132_1722 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1731_inst
    process(shl134_1727, conv107_1678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl134_1727, conv107_1678, tmp_var);
      add135_1732 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1736_inst
    process(add135_1732, conv98_1619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add135_1732, conv98_1619, tmp_var);
      add142_1737 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1741_inst
    process(add135_1732, conv100_1623) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add135_1732, conv100_1623, tmp_var);
      add146_1742 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1746_inst
    process(add101_1638, add135_1732) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add101_1638, add135_1732, tmp_var);
      add149_1747 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1559_inst
    process(iNsTr_14_1554) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_14_1554, type_cast_1558_wire_constant, tmp_var);
      xx_xop_1560 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1584_inst
    process(iNsTr_20_1570) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_20_1570, type_cast_1583_wire_constant, tmp_var);
      indvarx_xnext_1585 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1764_inst
    process(inc152_1760, shr79194_1606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc152_1760, shr79194_1606, tmp_var);
      cmp157_1765 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1788_inst
    process(inc160x_xcolx_x1_1777, add33_1444) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc160x_xcolx_x1_1777, add33_1444, tmp_var);
      cmp165_1789 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1812_inst
    process(inc169x_xrowx_x1_1801, add13_1394) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc169x_xrowx_x1_1801, add13_1394, tmp_var);
      cmp175_1813 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1589_inst
    process(indvarx_xnext_1585, tmp204_1567) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1585, tmp204_1567, tmp_var);
      exitcond1_1590 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1605_inst
    process(add53_1494) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add53_1494, type_cast_1604_wire_constant, tmp_var);
      shr79194_1606 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1537_inst
    process(tmp199_1532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp199_1532, type_cast_1536_wire_constant, tmp_var);
      tmp200_1538 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1610_inst
    process(shr79194_1606, add23_1419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(shr79194_1606, add23_1419, tmp_var);
      mul86_1611 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1503_inst
    process(conv59_1499, add_1369) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv59_1499, add_1369, tmp_var);
      mul_1504 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1508_inst
    process(mul_1504, add43_1469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1504, add43_1469, tmp_var);
      mul62_1509 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1526_inst
    process(add_1369, add43_1469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1369, add43_1469, tmp_var);
      tmp_1527 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1531_inst
    process(tmp_1527, conv59_1499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1527, conv59_1499, tmp_var);
      tmp199_1532 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1690_inst
    process(conv115_1686, conv113_1627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_1686, conv113_1627, tmp_var);
      mul116_1691 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1700_inst
    process(add117_1696, conv98_1619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add117_1696, conv98_1619, tmp_var);
      mul118_1701 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1716_inst
    process(conv115_1686, conv59_1499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_1686, conv59_1499, tmp_var);
      mul131_1717 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1726_inst
    process(mul133_1633, add132_1722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul133_1633, add132_1722, tmp_var);
      shl134_1727 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1859_inst
    process(conv113_1627, conv189_1851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv113_1627, conv189_1851, tmp_var);
      mul190_1860 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1864_inst
    process(mul190_1860, conv192_1855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul190_1860, conv192_1855, tmp_var);
      mul193_1865 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1819_inst
    process(cmp175_1813) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp175_1813, tmp_var);
      NOT_u1_u1_1819_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1393_inst
    process(shl10_1382, conv12_1389) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1382, conv12_1389, tmp_var);
      add13_1394 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1418_inst
    process(shl20_1407, conv22_1414) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1407, conv22_1414, tmp_var);
      add23_1419 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1443_inst
    process(shl30_1432, conv32_1439) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1432, conv32_1439, tmp_var);
      add33_1444 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1493_inst
    process(shl50_1482, conv52_1489) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1482, conv52_1489, tmp_var);
      add53_1494 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1368_inst
    process(shl_1357, conv3_1364) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1357, conv3_1364, tmp_var);
      add_1369 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1468_inst
    process(shl40_1457, conv42_1464) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1457, conv42_1464, tmp_var);
      add43_1469 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1381_inst
    process(conv9_1376) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1376, type_cast_1380_wire_constant, tmp_var);
      shl10_1382 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1406_inst
    process(conv19_1401) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1401, type_cast_1405_wire_constant, tmp_var);
      shl20_1407 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1431_inst
    process(conv29_1426) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1426, type_cast_1430_wire_constant, tmp_var);
      shl30_1432 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1481_inst
    process(conv49_1476) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1476, type_cast_1480_wire_constant, tmp_var);
      shl50_1482 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1356_inst
    process(conv1_1351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1351, type_cast_1355_wire_constant, tmp_var);
      shl_1357 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1456_inst
    process(conv39_1451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1451, type_cast_1455_wire_constant, tmp_var);
      shl40_1457 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1632_inst
    process(conv98_1619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_1619, type_cast_1631_wire_constant, tmp_var);
      mul133_1633 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1711_inst
    process(add119_1706) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add119_1706, type_cast_1710_wire_constant, tmp_var);
      shl120_1712 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1842_inst
    process(conv181_1838, conv90_1830) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv181_1838, conv90_1830, tmp_var);
      sub_1843 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1514_inst
    process(mul62_1509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul62_1509, type_cast_1513_wire_constant, tmp_var);
      cmp196_1515 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1543_inst
    process(tmp200_1538) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp200_1538, type_cast_1542_wire_constant, tmp_var);
      tmp201_1544 <= tmp_var; --
    end process;
    -- unary operator type_cast_1828_inst
    process(call89_1614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call89_1614, tmp_var);
      type_cast_1828_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1836_inst
    process(call180_1833) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call180_1833, tmp_var);
      type_cast_1836_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_1484_inst RPIPE_maxpool_input_pipe_1471_inst RPIPE_maxpool_input_pipe_1459_inst RPIPE_maxpool_input_pipe_1446_inst RPIPE_maxpool_input_pipe_1434_inst RPIPE_maxpool_input_pipe_1346_inst RPIPE_maxpool_input_pipe_1359_inst RPIPE_maxpool_input_pipe_1371_inst RPIPE_maxpool_input_pipe_1384_inst RPIPE_maxpool_input_pipe_1396_inst RPIPE_maxpool_input_pipe_1409_inst RPIPE_maxpool_input_pipe_1421_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(95 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1484_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1471_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1459_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1446_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1434_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1346_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1359_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1371_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1384_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1396_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1409_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1421_inst_req_0;
      RPIPE_maxpool_input_pipe_1484_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1471_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1459_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1446_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1434_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1346_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1359_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1371_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1384_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1396_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1409_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1421_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1484_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1471_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1459_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1446_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1434_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1346_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1359_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1371_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1384_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1396_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1409_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1421_inst_req_1;
      RPIPE_maxpool_input_pipe_1484_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1471_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1459_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1446_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1434_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1346_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1359_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1371_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1384_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1396_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1409_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1421_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call51_1485 <= data_out(95 downto 88);
      call46_1472 <= data_out(87 downto 80);
      call41_1460 <= data_out(79 downto 72);
      call36_1447 <= data_out(71 downto 64);
      call31_1435 <= data_out(63 downto 56);
      call_1347 <= data_out(55 downto 48);
      call2_1360 <= data_out(47 downto 40);
      call6_1372 <= data_out(39 downto 32);
      call11_1385 <= data_out(31 downto 24);
      call16_1397 <= data_out(23 downto 16);
      call21_1410 <= data_out(15 downto 8);
      call26_1422 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1844_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1844_inst_req_0;
      WPIPE_elapsed_time_pipe_1844_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1844_inst_req_1;
      WPIPE_elapsed_time_pipe_1844_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1843;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1579_call 
    fill_T_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1579_call_req_0;
      call_stmt_1579_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1579_call_req_1;
      call_stmt_1579_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_T_call_group_0_gI: SplitGuardInterface generic map(name => "fill_T_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_20_1570;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_T_call_reqs(0),
          ackR => fill_T_call_acks(0),
          dataR => fill_T_call_data(63 downto 0),
          tagR => fill_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_T_return_acks(0), -- cross-over
          ackL => fill_T_return_reqs(0), -- cross-over
          tagL => fill_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1833_call call_stmt_1614_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1833_call_req_0;
      reqL_unguarded(0) <= call_stmt_1614_call_req_0;
      call_stmt_1833_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1614_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1833_call_req_1;
      reqR_unguarded(0) <= call_stmt_1614_call_req_1;
      call_stmt_1833_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1614_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call180_1833 <= data_out(127 downto 64);
      call89_1614 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1754_call 
    maxPool4_call_group_2: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1754_call_req_0;
      call_stmt_1754_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1754_call_req_1;
      call_stmt_1754_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_2_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= shl120_1712 & add135_1732 & add142_1737 & add146_1742 & add149_1747;
      call150_1754 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 160,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(159 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1867_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1867_call_req_0;
      call_stmt_1867_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1867_call_req_1;
      call_stmt_1867_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul193_1865;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end maxPool3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    output : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 160)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_360_start: Boolean;
  signal maxPool4_CP_360_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u32_u64_1064_inst_ack_0 : boolean;
  signal slice_255_inst_ack_1 : boolean;
  signal slice_379_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1090_inst_req_0 : boolean;
  signal W_myptr5_1049_delayed_8_0_1049_inst_ack_0 : boolean;
  signal slice_275_inst_req_1 : boolean;
  signal slice_255_inst_req_1 : boolean;
  signal slice_247_inst_req_0 : boolean;
  signal slice_247_inst_ack_0 : boolean;
  signal W_myptr5_1049_delayed_8_0_1049_inst_ack_1 : boolean;
  signal slice_255_inst_ack_0 : boolean;
  signal slice_223_inst_ack_1 : boolean;
  signal slice_243_inst_ack_0 : boolean;
  signal slice_243_inst_req_0 : boolean;
  signal slice_251_inst_ack_0 : boolean;
  signal slice_255_inst_req_0 : boolean;
  signal slice_387_inst_req_0 : boolean;
  signal slice_263_inst_ack_0 : boolean;
  signal slice_223_inst_req_0 : boolean;
  signal slice_235_inst_ack_1 : boolean;
  signal slice_235_inst_req_1 : boolean;
  signal slice_239_inst_req_0 : boolean;
  signal W_myptr6_1072_delayed_8_0_1075_inst_ack_0 : boolean;
  signal ptr_deref_1053_store_0_req_1 : boolean;
  signal slice_223_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1064_inst_req_0 : boolean;
  signal slice_251_inst_req_0 : boolean;
  signal addr_of_1047_final_reg_req_0 : boolean;
  signal slice_259_inst_ack_1 : boolean;
  signal slice_235_inst_ack_0 : boolean;
  signal slice_259_inst_req_1 : boolean;
  signal slice_235_inst_req_0 : boolean;
  signal slice_243_inst_ack_1 : boolean;
  signal slice_223_inst_ack_0 : boolean;
  signal slice_271_inst_ack_0 : boolean;
  signal slice_267_inst_ack_1 : boolean;
  signal slice_259_inst_ack_0 : boolean;
  signal array_obj_ref_1072_index_offset_req_0 : boolean;
  signal slice_399_inst_ack_0 : boolean;
  signal slice_399_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1064_inst_req_1 : boolean;
  signal slice_251_inst_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_ack_0 : boolean;
  signal slice_379_inst_req_1 : boolean;
  signal slice_247_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1064_inst_ack_1 : boolean;
  signal slice_379_inst_ack_1 : boolean;
  signal slice_259_inst_req_0 : boolean;
  signal slice_231_inst_ack_1 : boolean;
  signal slice_231_inst_req_1 : boolean;
  signal slice_251_inst_req_1 : boolean;
  signal addr_of_1047_final_reg_ack_0 : boolean;
  signal slice_239_inst_ack_1 : boolean;
  signal array_obj_ref_1072_index_offset_req_1 : boolean;
  signal slice_231_inst_ack_0 : boolean;
  signal slice_231_inst_req_0 : boolean;
  signal slice_267_inst_req_1 : boolean;
  signal slice_275_inst_req_0 : boolean;
  signal slice_271_inst_ack_1 : boolean;
  signal slice_271_inst_req_1 : boolean;
  signal slice_379_inst_ack_0 : boolean;
  signal slice_247_inst_req_1 : boolean;
  signal slice_275_inst_ack_0 : boolean;
  signal slice_275_inst_ack_1 : boolean;
  signal slice_263_inst_ack_1 : boolean;
  signal slice_227_inst_ack_0 : boolean;
  signal slice_263_inst_req_1 : boolean;
  signal slice_227_inst_req_0 : boolean;
  signal W_myptr6_1072_delayed_8_0_1075_inst_req_0 : boolean;
  signal W_myptr5_1049_delayed_8_0_1049_inst_req_1 : boolean;
  signal slice_271_inst_req_0 : boolean;
  signal slice_263_inst_req_0 : boolean;
  signal slice_383_inst_req_0 : boolean;
  signal addr_of_126_final_reg_req_0 : boolean;
  signal addr_of_126_final_reg_ack_0 : boolean;
  signal slice_383_inst_ack_0 : boolean;
  signal addr_of_126_final_reg_req_1 : boolean;
  signal addr_of_126_final_reg_ack_1 : boolean;
  signal addr_of_1073_final_reg_ack_1 : boolean;
  signal slice_219_inst_ack_1 : boolean;
  signal slice_267_inst_ack_0 : boolean;
  signal slice_227_inst_ack_1 : boolean;
  signal slice_219_inst_req_1 : boolean;
  signal slice_399_inst_req_0 : boolean;
  signal slice_227_inst_req_1 : boolean;
  signal slice_267_inst_req_0 : boolean;
  signal ptr_deref_1053_store_0_ack_1 : boolean;
  signal CONCAT_u32_u64_1090_inst_ack_0 : boolean;
  signal slice_239_inst_req_1 : boolean;
  signal slice_243_inst_req_1 : boolean;
  signal slice_399_inst_req_1 : boolean;
  signal slice_239_inst_ack_0 : boolean;
  signal slice_219_inst_ack_0 : boolean;
  signal slice_219_inst_req_0 : boolean;
  signal array_obj_ref_1072_index_offset_ack_1 : boolean;
  signal slice_387_inst_ack_0 : boolean;
  signal addr_of_1047_final_reg_req_1 : boolean;
  signal slice_387_inst_req_1 : boolean;
  signal addr_of_1073_final_reg_req_0 : boolean;
  signal W_myptr6_1072_delayed_8_0_1075_inst_req_1 : boolean;
  signal array_obj_ref_104_index_offset_req_0 : boolean;
  signal array_obj_ref_104_index_offset_ack_0 : boolean;
  signal array_obj_ref_104_index_offset_req_1 : boolean;
  signal array_obj_ref_104_index_offset_ack_1 : boolean;
  signal W_myptr6_1072_delayed_8_0_1075_inst_ack_1 : boolean;
  signal addr_of_105_final_reg_req_0 : boolean;
  signal addr_of_105_final_reg_ack_0 : boolean;
  signal addr_of_105_final_reg_req_1 : boolean;
  signal addr_of_105_final_reg_ack_1 : boolean;
  signal slice_387_inst_ack_1 : boolean;
  signal addr_of_1073_final_reg_ack_0 : boolean;
  signal array_obj_ref_111_index_offset_req_0 : boolean;
  signal array_obj_ref_111_index_offset_ack_0 : boolean;
  signal array_obj_ref_111_index_offset_req_1 : boolean;
  signal array_obj_ref_111_index_offset_ack_1 : boolean;
  signal addr_of_1047_final_reg_ack_1 : boolean;
  signal addr_of_112_final_reg_req_0 : boolean;
  signal addr_of_112_final_reg_ack_0 : boolean;
  signal addr_of_112_final_reg_req_1 : boolean;
  signal addr_of_112_final_reg_ack_1 : boolean;
  signal array_obj_ref_118_index_offset_req_0 : boolean;
  signal array_obj_ref_118_index_offset_ack_0 : boolean;
  signal array_obj_ref_118_index_offset_req_1 : boolean;
  signal array_obj_ref_118_index_offset_ack_1 : boolean;
  signal addr_of_119_final_reg_req_0 : boolean;
  signal addr_of_119_final_reg_ack_0 : boolean;
  signal addr_of_119_final_reg_req_1 : boolean;
  signal addr_of_119_final_reg_ack_1 : boolean;
  signal addr_of_1073_final_reg_req_1 : boolean;
  signal array_obj_ref_125_index_offset_req_0 : boolean;
  signal array_obj_ref_125_index_offset_ack_0 : boolean;
  signal array_obj_ref_125_index_offset_req_1 : boolean;
  signal array_obj_ref_125_index_offset_ack_1 : boolean;
  signal ptr_deref_130_load_0_req_0 : boolean;
  signal ptr_deref_130_load_0_ack_0 : boolean;
  signal ptr_deref_130_load_0_req_1 : boolean;
  signal ptr_deref_130_load_0_ack_1 : boolean;
  signal array_obj_ref_1046_index_offset_req_0 : boolean;
  signal slice_383_inst_req_1 : boolean;
  signal ptr_deref_134_load_0_req_0 : boolean;
  signal ptr_deref_134_load_0_ack_0 : boolean;
  signal ptr_deref_134_load_0_req_1 : boolean;
  signal ptr_deref_134_load_0_ack_1 : boolean;
  signal array_obj_ref_1046_index_offset_ack_0 : boolean;
  signal ptr_deref_1053_store_0_req_0 : boolean;
  signal W_myptr5_1049_delayed_8_0_1049_inst_req_0 : boolean;
  signal ptr_deref_138_load_0_req_0 : boolean;
  signal ptr_deref_138_load_0_ack_0 : boolean;
  signal slice_383_inst_ack_1 : boolean;
  signal ptr_deref_138_load_0_req_1 : boolean;
  signal ptr_deref_138_load_0_ack_1 : boolean;
  signal array_obj_ref_1046_index_offset_req_1 : boolean;
  signal ptr_deref_142_load_0_req_0 : boolean;
  signal ptr_deref_142_load_0_ack_0 : boolean;
  signal ptr_deref_142_load_0_req_1 : boolean;
  signal ptr_deref_142_load_0_ack_1 : boolean;
  signal slice_147_inst_req_0 : boolean;
  signal slice_147_inst_ack_0 : boolean;
  signal slice_147_inst_req_1 : boolean;
  signal slice_147_inst_ack_1 : boolean;
  signal slice_151_inst_req_0 : boolean;
  signal slice_151_inst_ack_0 : boolean;
  signal slice_151_inst_req_1 : boolean;
  signal slice_151_inst_ack_1 : boolean;
  signal slice_155_inst_req_0 : boolean;
  signal slice_155_inst_ack_0 : boolean;
  signal slice_155_inst_req_1 : boolean;
  signal slice_155_inst_ack_1 : boolean;
  signal slice_159_inst_req_0 : boolean;
  signal slice_159_inst_ack_0 : boolean;
  signal slice_159_inst_req_1 : boolean;
  signal slice_159_inst_ack_1 : boolean;
  signal slice_163_inst_req_0 : boolean;
  signal slice_163_inst_ack_0 : boolean;
  signal slice_163_inst_req_1 : boolean;
  signal slice_163_inst_ack_1 : boolean;
  signal slice_167_inst_req_0 : boolean;
  signal slice_167_inst_ack_0 : boolean;
  signal slice_167_inst_req_1 : boolean;
  signal slice_167_inst_ack_1 : boolean;
  signal slice_171_inst_req_0 : boolean;
  signal slice_171_inst_ack_0 : boolean;
  signal slice_171_inst_req_1 : boolean;
  signal slice_171_inst_ack_1 : boolean;
  signal slice_175_inst_req_0 : boolean;
  signal slice_175_inst_ack_0 : boolean;
  signal slice_175_inst_req_1 : boolean;
  signal slice_175_inst_ack_1 : boolean;
  signal slice_179_inst_req_0 : boolean;
  signal slice_179_inst_ack_0 : boolean;
  signal slice_179_inst_req_1 : boolean;
  signal slice_179_inst_ack_1 : boolean;
  signal slice_183_inst_req_0 : boolean;
  signal slice_183_inst_ack_0 : boolean;
  signal slice_183_inst_req_1 : boolean;
  signal slice_183_inst_ack_1 : boolean;
  signal slice_187_inst_req_0 : boolean;
  signal slice_187_inst_ack_0 : boolean;
  signal slice_187_inst_req_1 : boolean;
  signal slice_187_inst_ack_1 : boolean;
  signal slice_191_inst_req_0 : boolean;
  signal slice_191_inst_ack_0 : boolean;
  signal slice_191_inst_req_1 : boolean;
  signal slice_191_inst_ack_1 : boolean;
  signal slice_195_inst_req_0 : boolean;
  signal slice_195_inst_ack_0 : boolean;
  signal slice_195_inst_req_1 : boolean;
  signal slice_195_inst_ack_1 : boolean;
  signal slice_199_inst_req_0 : boolean;
  signal slice_199_inst_ack_0 : boolean;
  signal slice_199_inst_req_1 : boolean;
  signal slice_199_inst_ack_1 : boolean;
  signal slice_203_inst_req_0 : boolean;
  signal slice_203_inst_ack_0 : boolean;
  signal slice_203_inst_req_1 : boolean;
  signal slice_203_inst_ack_1 : boolean;
  signal slice_207_inst_req_0 : boolean;
  signal slice_207_inst_ack_0 : boolean;
  signal slice_207_inst_req_1 : boolean;
  signal slice_207_inst_ack_1 : boolean;
  signal slice_211_inst_req_0 : boolean;
  signal slice_211_inst_ack_0 : boolean;
  signal slice_211_inst_req_1 : boolean;
  signal slice_211_inst_ack_1 : boolean;
  signal slice_215_inst_req_0 : boolean;
  signal slice_215_inst_ack_0 : boolean;
  signal slice_215_inst_req_1 : boolean;
  signal slice_215_inst_ack_1 : boolean;
  signal slice_395_inst_ack_1 : boolean;
  signal slice_279_inst_req_0 : boolean;
  signal slice_279_inst_ack_0 : boolean;
  signal slice_279_inst_req_1 : boolean;
  signal slice_279_inst_ack_1 : boolean;
  signal slice_395_inst_req_1 : boolean;
  signal array_obj_ref_1046_index_offset_ack_1 : boolean;
  signal slice_283_inst_req_0 : boolean;
  signal slice_283_inst_ack_0 : boolean;
  signal slice_283_inst_req_1 : boolean;
  signal slice_283_inst_ack_1 : boolean;
  signal slice_287_inst_req_0 : boolean;
  signal slice_287_inst_ack_0 : boolean;
  signal ptr_deref_1053_store_0_ack_0 : boolean;
  signal slice_287_inst_req_1 : boolean;
  signal slice_287_inst_ack_1 : boolean;
  signal slice_395_inst_ack_0 : boolean;
  signal slice_291_inst_req_0 : boolean;
  signal slice_291_inst_ack_0 : boolean;
  signal slice_395_inst_req_0 : boolean;
  signal slice_291_inst_req_1 : boolean;
  signal slice_291_inst_ack_1 : boolean;
  signal slice_295_inst_req_0 : boolean;
  signal slice_295_inst_ack_0 : boolean;
  signal slice_375_inst_ack_1 : boolean;
  signal slice_295_inst_req_1 : boolean;
  signal slice_295_inst_ack_1 : boolean;
  signal slice_375_inst_req_1 : boolean;
  signal slice_299_inst_req_0 : boolean;
  signal slice_299_inst_ack_0 : boolean;
  signal slice_299_inst_req_1 : boolean;
  signal slice_299_inst_ack_1 : boolean;
  signal slice_391_inst_ack_1 : boolean;
  signal slice_391_inst_req_1 : boolean;
  signal slice_375_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1090_inst_ack_1 : boolean;
  signal slice_375_inst_req_0 : boolean;
  signal slice_303_inst_req_0 : boolean;
  signal slice_303_inst_ack_0 : boolean;
  signal slice_303_inst_req_1 : boolean;
  signal slice_303_inst_ack_1 : boolean;
  signal slice_391_inst_ack_0 : boolean;
  signal slice_307_inst_req_0 : boolean;
  signal slice_307_inst_ack_0 : boolean;
  signal slice_307_inst_req_1 : boolean;
  signal slice_307_inst_ack_1 : boolean;
  signal slice_391_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1090_inst_req_1 : boolean;
  signal slice_311_inst_req_0 : boolean;
  signal slice_311_inst_ack_0 : boolean;
  signal slice_311_inst_req_1 : boolean;
  signal slice_311_inst_ack_1 : boolean;
  signal slice_315_inst_req_0 : boolean;
  signal slice_315_inst_ack_0 : boolean;
  signal slice_315_inst_req_1 : boolean;
  signal slice_315_inst_ack_1 : boolean;
  signal slice_319_inst_req_0 : boolean;
  signal slice_319_inst_ack_0 : boolean;
  signal slice_319_inst_req_1 : boolean;
  signal slice_319_inst_ack_1 : boolean;
  signal slice_323_inst_req_0 : boolean;
  signal slice_323_inst_ack_0 : boolean;
  signal slice_323_inst_req_1 : boolean;
  signal slice_323_inst_ack_1 : boolean;
  signal slice_327_inst_req_0 : boolean;
  signal slice_327_inst_ack_0 : boolean;
  signal slice_327_inst_req_1 : boolean;
  signal slice_327_inst_ack_1 : boolean;
  signal slice_331_inst_req_0 : boolean;
  signal slice_331_inst_ack_0 : boolean;
  signal slice_331_inst_req_1 : boolean;
  signal slice_331_inst_ack_1 : boolean;
  signal slice_335_inst_req_0 : boolean;
  signal slice_335_inst_ack_0 : boolean;
  signal slice_335_inst_req_1 : boolean;
  signal slice_335_inst_ack_1 : boolean;
  signal slice_339_inst_req_0 : boolean;
  signal slice_339_inst_ack_0 : boolean;
  signal slice_339_inst_req_1 : boolean;
  signal slice_339_inst_ack_1 : boolean;
  signal slice_343_inst_req_0 : boolean;
  signal slice_343_inst_ack_0 : boolean;
  signal slice_343_inst_req_1 : boolean;
  signal slice_343_inst_ack_1 : boolean;
  signal slice_347_inst_req_0 : boolean;
  signal slice_347_inst_ack_0 : boolean;
  signal slice_347_inst_req_1 : boolean;
  signal slice_347_inst_ack_1 : boolean;
  signal slice_351_inst_req_0 : boolean;
  signal slice_351_inst_ack_0 : boolean;
  signal slice_351_inst_req_1 : boolean;
  signal slice_351_inst_ack_1 : boolean;
  signal slice_355_inst_req_0 : boolean;
  signal slice_355_inst_ack_0 : boolean;
  signal slice_355_inst_req_1 : boolean;
  signal slice_355_inst_ack_1 : boolean;
  signal slice_359_inst_req_0 : boolean;
  signal slice_359_inst_ack_0 : boolean;
  signal slice_359_inst_req_1 : boolean;
  signal slice_359_inst_ack_1 : boolean;
  signal slice_363_inst_req_0 : boolean;
  signal slice_363_inst_ack_0 : boolean;
  signal slice_363_inst_req_1 : boolean;
  signal slice_363_inst_ack_1 : boolean;
  signal slice_367_inst_req_0 : boolean;
  signal slice_367_inst_ack_0 : boolean;
  signal slice_367_inst_req_1 : boolean;
  signal slice_367_inst_ack_1 : boolean;
  signal slice_371_inst_req_0 : boolean;
  signal slice_371_inst_ack_0 : boolean;
  signal slice_371_inst_req_1 : boolean;
  signal slice_371_inst_ack_1 : boolean;
  signal ptr_deref_1079_store_0_req_0 : boolean;
  signal ptr_deref_1079_store_0_ack_0 : boolean;
  signal ptr_deref_1079_store_0_req_1 : boolean;
  signal ptr_deref_1079_store_0_ack_1 : boolean;
  signal array_obj_ref_1098_index_offset_req_0 : boolean;
  signal array_obj_ref_1098_index_offset_ack_0 : boolean;
  signal array_obj_ref_1098_index_offset_req_1 : boolean;
  signal array_obj_ref_1098_index_offset_ack_1 : boolean;
  signal addr_of_1099_final_reg_req_0 : boolean;
  signal addr_of_1099_final_reg_ack_0 : boolean;
  signal addr_of_1099_final_reg_req_1 : boolean;
  signal addr_of_1099_final_reg_ack_1 : boolean;
  signal W_myptr7_1095_delayed_8_0_1101_inst_req_0 : boolean;
  signal W_myptr7_1095_delayed_8_0_1101_inst_ack_0 : boolean;
  signal W_myptr7_1095_delayed_8_0_1101_inst_req_1 : boolean;
  signal W_myptr7_1095_delayed_8_0_1101_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1116_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1116_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1116_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1116_inst_ack_1 : boolean;
  signal ptr_deref_1105_store_0_req_0 : boolean;
  signal ptr_deref_1105_store_0_ack_0 : boolean;
  signal ptr_deref_1105_store_0_req_1 : boolean;
  signal ptr_deref_1105_store_0_ack_1 : boolean;
  signal array_obj_ref_1124_index_offset_req_0 : boolean;
  signal array_obj_ref_1124_index_offset_ack_0 : boolean;
  signal array_obj_ref_1124_index_offset_req_1 : boolean;
  signal array_obj_ref_1124_index_offset_ack_1 : boolean;
  signal addr_of_1125_final_reg_req_0 : boolean;
  signal addr_of_1125_final_reg_ack_0 : boolean;
  signal addr_of_1125_final_reg_req_1 : boolean;
  signal addr_of_1125_final_reg_ack_1 : boolean;
  signal W_myptr8_1118_delayed_8_0_1127_inst_req_0 : boolean;
  signal W_myptr8_1118_delayed_8_0_1127_inst_ack_0 : boolean;
  signal W_myptr8_1118_delayed_8_0_1127_inst_req_1 : boolean;
  signal W_myptr8_1118_delayed_8_0_1127_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1142_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1142_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1142_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1142_inst_ack_1 : boolean;
  signal ptr_deref_1131_store_0_req_0 : boolean;
  signal ptr_deref_1131_store_0_ack_0 : boolean;
  signal ptr_deref_1131_store_0_req_1 : boolean;
  signal ptr_deref_1131_store_0_ack_1 : boolean;
  signal type_cast_1146_inst_req_0 : boolean;
  signal type_cast_1146_inst_ack_0 : boolean;
  signal type_cast_1146_inst_req_1 : boolean;
  signal type_cast_1146_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 160) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(tag_length + 159 downto 160) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 159 downto 160);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_360_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_360_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_360_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_360_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_360: Block -- control-path 
    signal maxPool4_CP_360_elements: BooleanArray(398 downto 0);
    -- 
  begin -- 
    maxPool4_CP_360_elements(0) <= maxPool4_CP_360_start;
    maxPool4_CP_360_symbol <= maxPool4_CP_360_elements(398);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	31 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	309 
    -- CP-element group 1: 	310 
    -- CP-element group 1: 	311 
    -- CP-element group 1: 	328 
    -- CP-element group 1: 	329 
    -- CP-element group 1: 	330 
    -- CP-element group 1: 	347 
    -- CP-element group 1: 	348 
    -- CP-element group 1: 	349 
    -- CP-element group 1: 	366 
    -- CP-element group 1: 	367 
    -- CP-element group 1: 	368 
    -- CP-element group 1:  members (105) 
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_resized_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_computed_1
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Sample/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_104_index_offset_req_0); -- 
    req_448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_111_index_offset_req_0); -- 
    req_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_118_index_offset_req_0); -- 
    req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_125_index_offset_req_0); -- 
    req_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_1046_index_offset_req_0); -- 
    req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_1072_index_offset_req_0); -- 
    req_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_1098_index_offset_req_0); -- 
    req_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(1), ack => array_obj_ref_1124_index_offset_req_0); -- 
    maxPool4_CP_360_elements(1) <= maxPool4_CP_360_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	311 
    -- CP-element group 2: 	330 
    -- CP-element group 2: 	349 
    -- CP-element group 2: 	368 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	392 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_1147/addr_update_enable
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_1147/addr_update_enable_out
      -- 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(311) & maxPool4_CP_360_elements(330) & maxPool4_CP_360_elements(349) & maxPool4_CP_360_elements(368);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	393 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_1147/addr1_update_enable
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_1147/addr1_update_enable_out
      -- 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(11);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	394 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_1147/addr2_update_enable
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_1147/addr2_update_enable_out
      -- 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(18);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	395 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_1147/addr3_update_enable
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_1147/addr3_update_enable_out
      -- 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(25);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	396 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_106_to_assign_stmt_1147/addr4_update_enable
      -- CP-element group 6: 	 assign_stmt_106_to_assign_stmt_1147/addr4_update_enable_out
      -- 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(32);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	397 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	385 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_106_to_assign_stmt_1147/output_update_enable
      -- CP-element group 7: 	 assign_stmt_106_to_assign_stmt_1147/output_update_enable_in
      -- 
    maxPool4_CP_360_elements(7) <= maxPool4_CP_360_elements(397);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_sample_start_
      -- CP-element group 8: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_request/$entry
      -- CP-element group 8: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_request/req
      -- 
    req_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(8), ack => addr_of_105_final_reg_req_0); -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(12) & maxPool4_CP_360_elements(13);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	38 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_update_start_
      -- CP-element group 9: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_complete/$entry
      -- CP-element group 9: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_complete/req
      -- 
    req_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(9), ack => addr_of_105_final_reg_req_1); -- 
    maxPool4_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(14) & maxPool4_CP_360_elements(38);
      gj_maxPool4_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_update_start
      -- CP-element group 10: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Update/$entry
      -- CP-element group 10: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Update/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(10), ack => array_obj_ref_104_index_offset_req_1); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(12) & maxPool4_CP_360_elements(13);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	391 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_sample_complete
      -- CP-element group 11: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Sample/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_104_index_offset_ack_0, ack => maxPool4_CP_360_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_offset_calculated
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Update/$exit
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_final_index_sum_regn_Update/ack
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_104_base_plus_offset/sum_rename_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_104_index_offset_ack_1, ack => maxPool4_CP_360_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_sample_completed_
      -- CP-element group 13: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_request/$exit
      -- CP-element group 13: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_request/ack
      -- 
    ack_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_105_final_reg_ack_0, ack => maxPool4_CP_360_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (19) 
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_address_calculated
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_word_address_calculated
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_root_address_calculated
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_address_resized
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_update_completed_
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_complete/$exit
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_105_complete/ack
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_addr_resize/$entry
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_addr_resize/$exit
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_plus_offset/$entry
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_plus_offset/$exit
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_word_addrgen/$entry
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_word_addrgen/$exit
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_word_addrgen/root_register_req
      -- CP-element group 14: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_word_addrgen/root_register_ack
      -- 
    ack_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_105_final_reg_ack_1, ack => maxPool4_CP_360_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_sample_start_
      -- CP-element group 15: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_request/$entry
      -- CP-element group 15: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_request/req
      -- 
    req_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(15), ack => addr_of_112_final_reg_req_0); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(19) & maxPool4_CP_360_elements(20);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	42 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_update_start_
      -- CP-element group 16: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_complete/$entry
      -- CP-element group 16: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_complete/req
      -- 
    req_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(16), ack => addr_of_112_final_reg_req_1); -- 
    maxPool4_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(21) & maxPool4_CP_360_elements(42);
      gj_maxPool4_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Update/req
      -- 
    req_453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(17), ack => array_obj_ref_111_index_offset_req_1); -- 
    maxPool4_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(19) & maxPool4_CP_360_elements(20);
      gj_maxPool4_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	391 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Sample/ack
      -- 
    ack_449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_111_index_offset_ack_0, ack => maxPool4_CP_360_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_root_address_calculated
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_offset_calculated
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_111_base_plus_offset/sum_rename_ack
      -- 
    ack_454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_111_index_offset_ack_1, ack => maxPool4_CP_360_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_sample_completed_
      -- CP-element group 20: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_request/$exit
      -- CP-element group 20: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_request/ack
      -- 
    ack_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_112_final_reg_ack_0, ack => maxPool4_CP_360_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	40 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_update_completed_
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_complete/$exit
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_112_complete/ack
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_address_resized
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_word_addrgen/root_register_ack
      -- 
    ack_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_112_final_reg_ack_1, ack => maxPool4_CP_360_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_sample_start_
      -- CP-element group 22: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_request/$entry
      -- CP-element group 22: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_request/req
      -- 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(22), ack => addr_of_119_final_reg_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(26) & maxPool4_CP_360_elements(27);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_update_start_
      -- CP-element group 23: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_complete/$entry
      -- CP-element group 23: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_complete/req
      -- 
    req_514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(23), ack => addr_of_119_final_reg_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(28) & maxPool4_CP_360_elements(46);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_update_start
      -- CP-element group 24: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Update/$entry
      -- CP-element group 24: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Update/req
      -- 
    req_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(24), ack => array_obj_ref_118_index_offset_req_1); -- 
    maxPool4_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(26) & maxPool4_CP_360_elements(27);
      gj_maxPool4_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	391 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_sample_complete
      -- CP-element group 25: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Sample/ack
      -- 
    ack_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_118_index_offset_ack_0, ack => maxPool4_CP_360_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (8) 
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_offset_calculated
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Update/$exit
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_final_index_sum_regn_Update/ack
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_118_base_plus_offset/sum_rename_ack
      -- 
    ack_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_118_index_offset_ack_1, ack => maxPool4_CP_360_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_sample_completed_
      -- CP-element group 27: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_request/$exit
      -- CP-element group 27: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_request/ack
      -- 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_119_final_reg_ack_0, ack => maxPool4_CP_360_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	44 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28:  members (19) 
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_update_completed_
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_complete/$exit
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_119_complete/ack
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_address_calculated
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_word_address_calculated
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_address_resized
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_addr_resize/$entry
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_addr_resize/$exit
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_addr_resize/base_resize_req
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_addr_resize/base_resize_ack
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_word_addrgen/$entry
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_word_addrgen/$exit
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_word_addrgen/root_register_req
      -- CP-element group 28: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_word_addrgen/root_register_ack
      -- 
    ack_515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_119_final_reg_ack_1, ack => maxPool4_CP_360_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_request/$entry
      -- CP-element group 29: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_request/req
      -- CP-element group 29: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_sample_start_
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(29), ack => addr_of_126_final_reg_req_0); -- 
    maxPool4_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(33) & maxPool4_CP_360_elements(34);
      gj_maxPool4_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	50 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_complete/$entry
      -- CP-element group 30: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_complete/req
      -- CP-element group 30: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_update_start_
      -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(30), ack => addr_of_126_final_reg_req_1); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(35) & maxPool4_CP_360_elements(50);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: 	34 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_update_start
      -- CP-element group 31: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Update/$entry
      -- CP-element group 31: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Update/req
      -- 
    req_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(31), ack => array_obj_ref_125_index_offset_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(33) & maxPool4_CP_360_elements(34);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	1 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	391 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Sample/ack
      -- 
    ack_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_offset_ack_0, ack => maxPool4_CP_360_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (8) 
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_base_plus_offset/$entry
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_base_plus_offset/$exit
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_root_address_calculated
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_offset_calculated
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_125_final_index_sum_regn_Update/ack
      -- 
    ack_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_125_index_offset_ack_1, ack => maxPool4_CP_360_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_request/$exit
      -- CP-element group 34: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_request/ack
      -- CP-element group 34: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_sample_completed_
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_126_final_reg_ack_0, ack => maxPool4_CP_360_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	48 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	30 
    -- CP-element group 35:  members (19) 
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_complete/$exit
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_complete/ack
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_root_address_calculated
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_126_update_completed_
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_address_calculated
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_word_address_calculated
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_address_resized
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_addr_resize/$entry
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_addr_resize/$exit
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_plus_offset/$entry
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_plus_offset/$exit
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_word_addrgen/$entry
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_word_addrgen/$exit
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_word_addrgen/root_register_req
      -- CP-element group 35: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_word_addrgen/root_register_ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_126_final_reg_ack_1, ack => maxPool4_CP_360_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_sample_start_
      -- CP-element group 36: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/$entry
      -- CP-element group 36: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/word_0/rr
      -- 
    rr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(36), ack => ptr_deref_130_load_0_req_0); -- 
    maxPool4_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(14) & maxPool4_CP_360_elements(38);
      gj_maxPool4_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	74 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	94 
    -- CP-element group 37: 	98 
    -- CP-element group 37: 	102 
    -- CP-element group 37: 	106 
    -- CP-element group 37: 	110 
    -- CP-element group 37: 	114 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_update_start_
      -- CP-element group 37: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/$entry
      -- CP-element group 37: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/$entry
      -- CP-element group 37: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/word_0/cr
      -- 
    cr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(37), ack => ptr_deref_130_load_0_req_1); -- 
    maxPool4_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(54) & maxPool4_CP_360_elements(58) & maxPool4_CP_360_elements(62) & maxPool4_CP_360_elements(66) & maxPool4_CP_360_elements(70) & maxPool4_CP_360_elements(74) & maxPool4_CP_360_elements(78) & maxPool4_CP_360_elements(82) & maxPool4_CP_360_elements(86) & maxPool4_CP_360_elements(90) & maxPool4_CP_360_elements(94) & maxPool4_CP_360_elements(98) & maxPool4_CP_360_elements(102) & maxPool4_CP_360_elements(106) & maxPool4_CP_360_elements(110) & maxPool4_CP_360_elements(114);
      gj_maxPool4_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_sample_completed_
      -- CP-element group 38: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/$exit
      -- CP-element group 38: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Sample/word_access_start/word_0/ra
      -- 
    ra_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_130_load_0_ack_0, ack => maxPool4_CP_360_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	72 
    -- CP-element group 39: 	76 
    -- CP-element group 39: 	80 
    -- CP-element group 39: 	84 
    -- CP-element group 39: 	88 
    -- CP-element group 39: 	92 
    -- CP-element group 39: 	96 
    -- CP-element group 39: 	100 
    -- CP-element group 39: 	104 
    -- CP-element group 39: 	108 
    -- CP-element group 39: 	112 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_update_completed_
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/$exit
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/$exit
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/ptr_deref_130_Merge/$entry
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/ptr_deref_130_Merge/$exit
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/ptr_deref_130_Merge/merge_req
      -- CP-element group 39: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_130_Update/ptr_deref_130_Merge/merge_ack
      -- 
    ca_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_130_load_0_ack_1, ack => maxPool4_CP_360_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_sample_start_
      -- CP-element group 40: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/word_0/rr
      -- 
    rr_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(40), ack => ptr_deref_134_load_0_req_0); -- 
    maxPool4_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(21) & maxPool4_CP_360_elements(42);
      gj_maxPool4_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	118 
    -- CP-element group 41: 	122 
    -- CP-element group 41: 	126 
    -- CP-element group 41: 	130 
    -- CP-element group 41: 	134 
    -- CP-element group 41: 	138 
    -- CP-element group 41: 	142 
    -- CP-element group 41: 	146 
    -- CP-element group 41: 	150 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	158 
    -- CP-element group 41: 	162 
    -- CP-element group 41: 	166 
    -- CP-element group 41: 	170 
    -- CP-element group 41: 	174 
    -- CP-element group 41: 	178 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_update_start_
      -- CP-element group 41: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/$entry
      -- CP-element group 41: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/$entry
      -- CP-element group 41: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/word_0/cr
      -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(41), ack => ptr_deref_134_load_0_req_1); -- 
    maxPool4_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(118) & maxPool4_CP_360_elements(122) & maxPool4_CP_360_elements(126) & maxPool4_CP_360_elements(130) & maxPool4_CP_360_elements(134) & maxPool4_CP_360_elements(138) & maxPool4_CP_360_elements(142) & maxPool4_CP_360_elements(146) & maxPool4_CP_360_elements(150) & maxPool4_CP_360_elements(154) & maxPool4_CP_360_elements(158) & maxPool4_CP_360_elements(162) & maxPool4_CP_360_elements(166) & maxPool4_CP_360_elements(170) & maxPool4_CP_360_elements(174) & maxPool4_CP_360_elements(178);
      gj_maxPool4_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	16 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_sample_completed_
      -- CP-element group 42: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Sample/word_access_start/word_0/ra
      -- 
    ra_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_134_load_0_ack_0, ack => maxPool4_CP_360_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	116 
    -- CP-element group 43: 	120 
    -- CP-element group 43: 	124 
    -- CP-element group 43: 	128 
    -- CP-element group 43: 	132 
    -- CP-element group 43: 	136 
    -- CP-element group 43: 	140 
    -- CP-element group 43: 	144 
    -- CP-element group 43: 	148 
    -- CP-element group 43: 	152 
    -- CP-element group 43: 	156 
    -- CP-element group 43: 	160 
    -- CP-element group 43: 	164 
    -- CP-element group 43: 	168 
    -- CP-element group 43: 	172 
    -- CP-element group 43: 	176 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_update_completed_
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/$exit
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/ptr_deref_134_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/ptr_deref_134_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/ptr_deref_134_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_134_Update/ptr_deref_134_Merge/merge_ack
      -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_134_load_0_ack_1, ack => maxPool4_CP_360_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	28 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_sample_start_
      -- CP-element group 44: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/$entry
      -- CP-element group 44: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/$entry
      -- CP-element group 44: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/word_0/rr
      -- 
    rr_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(44), ack => ptr_deref_138_load_0_req_0); -- 
    maxPool4_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(28) & maxPool4_CP_360_elements(46);
      gj_maxPool4_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	182 
    -- CP-element group 45: 	186 
    -- CP-element group 45: 	190 
    -- CP-element group 45: 	194 
    -- CP-element group 45: 	198 
    -- CP-element group 45: 	202 
    -- CP-element group 45: 	206 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	214 
    -- CP-element group 45: 	218 
    -- CP-element group 45: 	222 
    -- CP-element group 45: 	226 
    -- CP-element group 45: 	230 
    -- CP-element group 45: 	234 
    -- CP-element group 45: 	238 
    -- CP-element group 45: 	242 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_update_start_
      -- CP-element group 45: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/$entry
      -- CP-element group 45: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/$entry
      -- CP-element group 45: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/word_0/cr
      -- 
    cr_705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(45), ack => ptr_deref_138_load_0_req_1); -- 
    maxPool4_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(182) & maxPool4_CP_360_elements(186) & maxPool4_CP_360_elements(190) & maxPool4_CP_360_elements(194) & maxPool4_CP_360_elements(198) & maxPool4_CP_360_elements(202) & maxPool4_CP_360_elements(206) & maxPool4_CP_360_elements(210) & maxPool4_CP_360_elements(214) & maxPool4_CP_360_elements(218) & maxPool4_CP_360_elements(222) & maxPool4_CP_360_elements(226) & maxPool4_CP_360_elements(230) & maxPool4_CP_360_elements(234) & maxPool4_CP_360_elements(238) & maxPool4_CP_360_elements(242);
      gj_maxPool4_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_sample_completed_
      -- CP-element group 46: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Sample/word_access_start/word_0/ra
      -- 
    ra_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_0, ack => maxPool4_CP_360_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	204 
    -- CP-element group 47: 	208 
    -- CP-element group 47: 	212 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	220 
    -- CP-element group 47: 	224 
    -- CP-element group 47: 	228 
    -- CP-element group 47: 	232 
    -- CP-element group 47: 	236 
    -- CP-element group 47: 	240 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_update_completed_
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/$exit
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/ptr_deref_138_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/ptr_deref_138_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/ptr_deref_138_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_138_Update/ptr_deref_138_Merge/merge_ack
      -- 
    ca_706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_1, ack => maxPool4_CP_360_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_sample_start_
      -- CP-element group 48: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/word_0/rr
      -- 
    rr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(48), ack => ptr_deref_142_load_0_req_0); -- 
    maxPool4_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(35) & maxPool4_CP_360_elements(50);
      gj_maxPool4_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	246 
    -- CP-element group 49: 	250 
    -- CP-element group 49: 	254 
    -- CP-element group 49: 	258 
    -- CP-element group 49: 	262 
    -- CP-element group 49: 	266 
    -- CP-element group 49: 	270 
    -- CP-element group 49: 	274 
    -- CP-element group 49: 	278 
    -- CP-element group 49: 	282 
    -- CP-element group 49: 	286 
    -- CP-element group 49: 	290 
    -- CP-element group 49: 	294 
    -- CP-element group 49: 	298 
    -- CP-element group 49: 	302 
    -- CP-element group 49: 	306 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_update_start_
      -- CP-element group 49: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/$entry
      -- CP-element group 49: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/$entry
      -- CP-element group 49: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/word_0/cr
      -- 
    cr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(49), ack => ptr_deref_142_load_0_req_1); -- 
    maxPool4_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(246) & maxPool4_CP_360_elements(250) & maxPool4_CP_360_elements(254) & maxPool4_CP_360_elements(258) & maxPool4_CP_360_elements(262) & maxPool4_CP_360_elements(266) & maxPool4_CP_360_elements(270) & maxPool4_CP_360_elements(274) & maxPool4_CP_360_elements(278) & maxPool4_CP_360_elements(282) & maxPool4_CP_360_elements(286) & maxPool4_CP_360_elements(290) & maxPool4_CP_360_elements(294) & maxPool4_CP_360_elements(298) & maxPool4_CP_360_elements(302) & maxPool4_CP_360_elements(306);
      gj_maxPool4_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	30 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_sample_completed_
      -- CP-element group 50: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Sample/word_access_start/word_0/ra
      -- 
    ra_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_142_load_0_ack_0, ack => maxPool4_CP_360_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	244 
    -- CP-element group 51: 	248 
    -- CP-element group 51: 	252 
    -- CP-element group 51: 	256 
    -- CP-element group 51: 	260 
    -- CP-element group 51: 	264 
    -- CP-element group 51: 	268 
    -- CP-element group 51: 	272 
    -- CP-element group 51: 	276 
    -- CP-element group 51: 	280 
    -- CP-element group 51: 	284 
    -- CP-element group 51: 	288 
    -- CP-element group 51: 	292 
    -- CP-element group 51: 	296 
    -- CP-element group 51: 	300 
    -- CP-element group 51: 	304 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_update_completed_
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/$exit
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/ptr_deref_142_Merge/$entry
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/ptr_deref_142_Merge/$exit
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/ptr_deref_142_Merge/merge_req
      -- CP-element group 51: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_142_Update/ptr_deref_142_Merge/merge_ack
      -- 
    ca_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_142_load_0_ack_1, ack => maxPool4_CP_360_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_sample_start_
      -- CP-element group 52: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Sample/rr
      -- 
    rr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(52), ack => slice_147_inst_req_0); -- 
    maxPool4_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(54);
      gj_maxPool4_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	321 
    -- CP-element group 53: 	386 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_update_start_
      -- CP-element group 53: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Update/$entry
      -- CP-element group 53: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Update/cr
      -- 
    cr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(53), ack => slice_147_inst_req_1); -- 
    maxPool4_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(55) & maxPool4_CP_360_elements(321) & maxPool4_CP_360_elements(386);
      gj_maxPool4_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_sample_completed_
      -- CP-element group 54: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Sample/ra
      -- 
    ra_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_0, ack => maxPool4_CP_360_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	319 
    -- CP-element group 55: 	384 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_update_completed_
      -- CP-element group 55: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Update/$exit
      -- CP-element group 55: 	 assign_stmt_106_to_assign_stmt_1147/slice_147_Update/ca
      -- 
    ca_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_1, ack => maxPool4_CP_360_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_sample_start_
      -- CP-element group 56: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Sample/rr
      -- 
    rr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(56), ack => slice_151_inst_req_0); -- 
    maxPool4_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(58);
      gj_maxPool4_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	321 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_update_start_
      -- CP-element group 57: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Update/$entry
      -- CP-element group 57: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Update/cr
      -- 
    cr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(57), ack => slice_151_inst_req_1); -- 
    maxPool4_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(59) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_sample_completed_
      -- CP-element group 58: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Sample/ra
      -- 
    ra_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_0, ack => maxPool4_CP_360_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	319 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_update_completed_
      -- CP-element group 59: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Update/$exit
      -- CP-element group 59: 	 assign_stmt_106_to_assign_stmt_1147/slice_151_Update/ca
      -- 
    ca_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_1, ack => maxPool4_CP_360_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_sample_start_
      -- CP-element group 60: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Sample/rr
      -- 
    rr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(60), ack => slice_155_inst_req_0); -- 
    maxPool4_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(62);
      gj_maxPool4_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	321 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_update_start_
      -- CP-element group 61: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Update/$entry
      -- CP-element group 61: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Update/cr
      -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(61), ack => slice_155_inst_req_1); -- 
    maxPool4_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(63) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_sample_completed_
      -- CP-element group 62: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Sample/ra
      -- 
    ra_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_0, ack => maxPool4_CP_360_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	319 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_update_completed_
      -- CP-element group 63: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Update/$exit
      -- CP-element group 63: 	 assign_stmt_106_to_assign_stmt_1147/slice_155_Update/ca
      -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_1, ack => maxPool4_CP_360_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_sample_start_
      -- CP-element group 64: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Sample/rr
      -- 
    rr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(64), ack => slice_159_inst_req_0); -- 
    maxPool4_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(66);
      gj_maxPool4_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	321 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_update_start_
      -- CP-element group 65: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Update/$entry
      -- CP-element group 65: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Update/cr
      -- 
    cr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(65), ack => slice_159_inst_req_1); -- 
    maxPool4_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(67) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_sample_completed_
      -- CP-element group 66: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Sample/ra
      -- 
    ra_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_159_inst_ack_0, ack => maxPool4_CP_360_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	319 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_update_completed_
      -- CP-element group 67: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Update/$exit
      -- CP-element group 67: 	 assign_stmt_106_to_assign_stmt_1147/slice_159_Update/ca
      -- 
    ca_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_159_inst_ack_1, ack => maxPool4_CP_360_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_sample_start_
      -- CP-element group 68: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Sample/$entry
      -- CP-element group 68: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Sample/rr
      -- 
    rr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(68), ack => slice_163_inst_req_0); -- 
    maxPool4_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(70);
      gj_maxPool4_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	340 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_update_start_
      -- CP-element group 69: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Update/$entry
      -- CP-element group 69: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Update/cr
      -- 
    cr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(69), ack => slice_163_inst_req_1); -- 
    maxPool4_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(71) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_sample_completed_
      -- CP-element group 70: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Sample/$exit
      -- CP-element group 70: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Sample/ra
      -- 
    ra_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_163_inst_ack_0, ack => maxPool4_CP_360_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	338 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_update_completed_
      -- CP-element group 71: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Update/$exit
      -- CP-element group 71: 	 assign_stmt_106_to_assign_stmt_1147/slice_163_Update/ca
      -- 
    ca_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_163_inst_ack_1, ack => maxPool4_CP_360_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	39 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_sample_start_
      -- CP-element group 72: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Sample/rr
      -- 
    rr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(72), ack => slice_167_inst_req_0); -- 
    maxPool4_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(74);
      gj_maxPool4_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	340 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_update_start_
      -- CP-element group 73: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Update/$entry
      -- CP-element group 73: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Update/cr
      -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(73), ack => slice_167_inst_req_1); -- 
    maxPool4_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(75) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	37 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_sample_completed_
      -- CP-element group 74: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Sample/ra
      -- 
    ra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_167_inst_ack_0, ack => maxPool4_CP_360_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	338 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_update_completed_
      -- CP-element group 75: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Update/$exit
      -- CP-element group 75: 	 assign_stmt_106_to_assign_stmt_1147/slice_167_Update/ca
      -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_167_inst_ack_1, ack => maxPool4_CP_360_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	39 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_sample_start_
      -- CP-element group 76: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Sample/rr
      -- 
    rr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(76), ack => slice_171_inst_req_0); -- 
    maxPool4_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(78);
      gj_maxPool4_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	340 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_update_start_
      -- CP-element group 77: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Update/$entry
      -- CP-element group 77: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Update/cr
      -- 
    cr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(77), ack => slice_171_inst_req_1); -- 
    maxPool4_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(79) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_sample_completed_
      -- CP-element group 78: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Sample/ra
      -- 
    ra_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_171_inst_ack_0, ack => maxPool4_CP_360_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	338 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_update_completed_
      -- CP-element group 79: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Update/$exit
      -- CP-element group 79: 	 assign_stmt_106_to_assign_stmt_1147/slice_171_Update/ca
      -- 
    ca_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_171_inst_ack_1, ack => maxPool4_CP_360_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	39 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_sample_start_
      -- CP-element group 80: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Sample/$entry
      -- CP-element group 80: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Sample/rr
      -- 
    rr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(80), ack => slice_175_inst_req_0); -- 
    maxPool4_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(82);
      gj_maxPool4_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	340 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_update_start_
      -- CP-element group 81: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Update/$entry
      -- CP-element group 81: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Update/cr
      -- 
    cr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(81), ack => slice_175_inst_req_1); -- 
    maxPool4_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(83) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_sample_completed_
      -- CP-element group 82: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Sample/ra
      -- 
    ra_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_175_inst_ack_0, ack => maxPool4_CP_360_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	338 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_update_completed_
      -- CP-element group 83: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Update/$exit
      -- CP-element group 83: 	 assign_stmt_106_to_assign_stmt_1147/slice_175_Update/ca
      -- 
    ca_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_175_inst_ack_1, ack => maxPool4_CP_360_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	39 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_sample_start_
      -- CP-element group 84: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Sample/$entry
      -- CP-element group 84: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Sample/rr
      -- 
    rr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(84), ack => slice_179_inst_req_0); -- 
    maxPool4_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(86);
      gj_maxPool4_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	359 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_update_start_
      -- CP-element group 85: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Update/$entry
      -- CP-element group 85: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Update/cr
      -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(85), ack => slice_179_inst_req_1); -- 
    maxPool4_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(87) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_sample_completed_
      -- CP-element group 86: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Sample/ra
      -- 
    ra_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_179_inst_ack_0, ack => maxPool4_CP_360_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	357 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_update_completed_
      -- CP-element group 87: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Update/$exit
      -- CP-element group 87: 	 assign_stmt_106_to_assign_stmt_1147/slice_179_Update/ca
      -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_179_inst_ack_1, ack => maxPool4_CP_360_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	39 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_sample_start_
      -- CP-element group 88: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Sample/rr
      -- 
    rr_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(88), ack => slice_183_inst_req_0); -- 
    maxPool4_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(90);
      gj_maxPool4_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	359 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_update_start_
      -- CP-element group 89: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Update/$entry
      -- CP-element group 89: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Update/cr
      -- 
    cr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(89), ack => slice_183_inst_req_1); -- 
    maxPool4_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(91) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_sample_completed_
      -- CP-element group 90: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Sample/$exit
      -- CP-element group 90: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Sample/ra
      -- 
    ra_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_183_inst_ack_0, ack => maxPool4_CP_360_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	357 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_update_completed_
      -- CP-element group 91: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Update/$exit
      -- CP-element group 91: 	 assign_stmt_106_to_assign_stmt_1147/slice_183_Update/ca
      -- 
    ca_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_183_inst_ack_1, ack => maxPool4_CP_360_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	39 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_sample_start_
      -- CP-element group 92: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Sample/rr
      -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(92), ack => slice_187_inst_req_0); -- 
    maxPool4_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(94);
      gj_maxPool4_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	359 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_update_start_
      -- CP-element group 93: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Update/$entry
      -- CP-element group 93: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Update/cr
      -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(93), ack => slice_187_inst_req_1); -- 
    maxPool4_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(95) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_sample_completed_
      -- CP-element group 94: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Sample/ra
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_187_inst_ack_0, ack => maxPool4_CP_360_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	357 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_update_completed_
      -- CP-element group 95: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Update/$exit
      -- CP-element group 95: 	 assign_stmt_106_to_assign_stmt_1147/slice_187_Update/ca
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_187_inst_ack_1, ack => maxPool4_CP_360_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	39 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_sample_start_
      -- CP-element group 96: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Sample/$entry
      -- CP-element group 96: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Sample/rr
      -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(96), ack => slice_191_inst_req_0); -- 
    maxPool4_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(98);
      gj_maxPool4_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	359 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_update_start_
      -- CP-element group 97: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Update/$entry
      -- CP-element group 97: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Update/cr
      -- 
    cr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(97), ack => slice_191_inst_req_1); -- 
    maxPool4_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(99) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	37 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_sample_completed_
      -- CP-element group 98: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Sample/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_191_inst_ack_0, ack => maxPool4_CP_360_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	357 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_update_completed_
      -- CP-element group 99: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Update/$exit
      -- CP-element group 99: 	 assign_stmt_106_to_assign_stmt_1147/slice_191_Update/ca
      -- 
    ca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_191_inst_ack_1, ack => maxPool4_CP_360_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	39 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_sample_start_
      -- CP-element group 100: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Sample/$entry
      -- CP-element group 100: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Sample/rr
      -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(100), ack => slice_195_inst_req_0); -- 
    maxPool4_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(102);
      gj_maxPool4_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	378 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_update_start_
      -- CP-element group 101: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Update/$entry
      -- CP-element group 101: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Update/cr
      -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(101), ack => slice_195_inst_req_1); -- 
    maxPool4_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(103) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_sample_completed_
      -- CP-element group 102: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Sample/ra
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_195_inst_ack_0, ack => maxPool4_CP_360_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	376 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_update_completed_
      -- CP-element group 103: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Update/$exit
      -- CP-element group 103: 	 assign_stmt_106_to_assign_stmt_1147/slice_195_Update/ca
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_195_inst_ack_1, ack => maxPool4_CP_360_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	39 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_sample_start_
      -- CP-element group 104: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Sample/$entry
      -- CP-element group 104: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Sample/rr
      -- 
    rr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(104), ack => slice_199_inst_req_0); -- 
    maxPool4_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(106);
      gj_maxPool4_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	378 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_update_start_
      -- CP-element group 105: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Update/$entry
      -- CP-element group 105: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Update/cr
      -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(105), ack => slice_199_inst_req_1); -- 
    maxPool4_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(107) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	37 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_sample_completed_
      -- CP-element group 106: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Sample/$exit
      -- CP-element group 106: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Sample/ra
      -- 
    ra_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_199_inst_ack_0, ack => maxPool4_CP_360_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	376 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_update_completed_
      -- CP-element group 107: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Update/$exit
      -- CP-element group 107: 	 assign_stmt_106_to_assign_stmt_1147/slice_199_Update/ca
      -- 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_199_inst_ack_1, ack => maxPool4_CP_360_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	39 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_sample_start_
      -- CP-element group 108: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Sample/rr
      -- 
    rr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(108), ack => slice_203_inst_req_0); -- 
    maxPool4_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(110);
      gj_maxPool4_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	378 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_update_start_
      -- CP-element group 109: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Update/$entry
      -- CP-element group 109: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Update/cr
      -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(109), ack => slice_203_inst_req_1); -- 
    maxPool4_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(111) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	37 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_sample_completed_
      -- CP-element group 110: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Sample/ra
      -- 
    ra_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_203_inst_ack_0, ack => maxPool4_CP_360_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	376 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_update_completed_
      -- CP-element group 111: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Update/$exit
      -- CP-element group 111: 	 assign_stmt_106_to_assign_stmt_1147/slice_203_Update/ca
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_203_inst_ack_1, ack => maxPool4_CP_360_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	39 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_sample_start_
      -- CP-element group 112: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Sample/$entry
      -- CP-element group 112: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Sample/rr
      -- 
    rr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(112), ack => slice_207_inst_req_0); -- 
    maxPool4_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(39) & maxPool4_CP_360_elements(114);
      gj_maxPool4_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	378 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_update_start_
      -- CP-element group 113: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Update/$entry
      -- CP-element group 113: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Update/cr
      -- 
    cr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(113), ack => slice_207_inst_req_1); -- 
    maxPool4_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(115) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	37 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_sample_completed_
      -- CP-element group 114: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Sample/$exit
      -- CP-element group 114: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Sample/ra
      -- 
    ra_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_207_inst_ack_0, ack => maxPool4_CP_360_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	376 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_update_completed_
      -- CP-element group 115: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Update/$exit
      -- CP-element group 115: 	 assign_stmt_106_to_assign_stmt_1147/slice_207_Update/ca
      -- 
    ca_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_207_inst_ack_1, ack => maxPool4_CP_360_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	43 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_sample_start_
      -- CP-element group 116: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Sample/$entry
      -- CP-element group 116: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Sample/rr
      -- 
    rr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(116), ack => slice_211_inst_req_0); -- 
    maxPool4_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(118);
      gj_maxPool4_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	321 
    -- CP-element group 117: 	386 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_update_start_
      -- CP-element group 117: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Update/$entry
      -- CP-element group 117: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Update/cr
      -- 
    cr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(117), ack => slice_211_inst_req_1); -- 
    maxPool4_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(119) & maxPool4_CP_360_elements(321) & maxPool4_CP_360_elements(386);
      gj_maxPool4_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	41 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_sample_completed_
      -- CP-element group 118: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Sample/ra
      -- 
    ra_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_211_inst_ack_0, ack => maxPool4_CP_360_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	319 
    -- CP-element group 119: 	384 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_update_completed_
      -- CP-element group 119: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Update/$exit
      -- CP-element group 119: 	 assign_stmt_106_to_assign_stmt_1147/slice_211_Update/ca
      -- 
    ca_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_211_inst_ack_1, ack => maxPool4_CP_360_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	43 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_sample_start_
      -- CP-element group 120: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Sample/$entry
      -- CP-element group 120: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Sample/rr
      -- 
    rr_1007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(120), ack => slice_215_inst_req_0); -- 
    maxPool4_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(122);
      gj_maxPool4_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	321 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_update_start_
      -- CP-element group 121: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Update/$entry
      -- CP-element group 121: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Update/cr
      -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(121), ack => slice_215_inst_req_1); -- 
    maxPool4_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(123) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	41 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_sample_completed_
      -- CP-element group 122: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Sample/ra
      -- 
    ra_1008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_215_inst_ack_0, ack => maxPool4_CP_360_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	319 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_update_completed_
      -- CP-element group 123: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Update/$exit
      -- CP-element group 123: 	 assign_stmt_106_to_assign_stmt_1147/slice_215_Update/ca
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_215_inst_ack_1, ack => maxPool4_CP_360_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	43 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Sample/rr
      -- CP-element group 124: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_sample_start_
      -- CP-element group 124: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Sample/$entry
      -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(124), ack => slice_219_inst_req_0); -- 
    maxPool4_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(126);
      gj_maxPool4_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	321 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Update/cr
      -- CP-element group 125: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Update/$entry
      -- CP-element group 125: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_update_start_
      -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(125), ack => slice_219_inst_req_1); -- 
    maxPool4_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(127) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	41 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Sample/ra
      -- CP-element group 126: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_sample_completed_
      -- CP-element group 126: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Sample/$exit
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_219_inst_ack_0, ack => maxPool4_CP_360_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	319 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Update/ca
      -- CP-element group 127: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_Update/$exit
      -- CP-element group 127: 	 assign_stmt_106_to_assign_stmt_1147/slice_219_update_completed_
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_219_inst_ack_1, ack => maxPool4_CP_360_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	43 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Sample/rr
      -- CP-element group 128: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Sample/$entry
      -- CP-element group 128: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_sample_start_
      -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(128), ack => slice_223_inst_req_0); -- 
    maxPool4_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(130);
      gj_maxPool4_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	321 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Update/cr
      -- CP-element group 129: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Update/$entry
      -- CP-element group 129: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_update_start_
      -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(129), ack => slice_223_inst_req_1); -- 
    maxPool4_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(131) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	41 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Sample/ra
      -- CP-element group 130: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Sample/$exit
      -- CP-element group 130: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_sample_completed_
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_223_inst_ack_0, ack => maxPool4_CP_360_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	319 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Update/ca
      -- CP-element group 131: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_Update/$exit
      -- CP-element group 131: 	 assign_stmt_106_to_assign_stmt_1147/slice_223_update_completed_
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_223_inst_ack_1, ack => maxPool4_CP_360_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	43 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Sample/rr
      -- CP-element group 132: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Sample/$entry
      -- CP-element group 132: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_sample_start_
      -- 
    rr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(132), ack => slice_227_inst_req_0); -- 
    maxPool4_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(134);
      gj_maxPool4_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	340 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Update/$entry
      -- CP-element group 133: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Update/cr
      -- CP-element group 133: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_update_start_
      -- 
    cr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(133), ack => slice_227_inst_req_1); -- 
    maxPool4_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(135) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	41 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Sample/ra
      -- CP-element group 134: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_sample_completed_
      -- 
    ra_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_227_inst_ack_0, ack => maxPool4_CP_360_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	338 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Update/$exit
      -- CP-element group 135: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_update_completed_
      -- CP-element group 135: 	 assign_stmt_106_to_assign_stmt_1147/slice_227_Update/ca
      -- 
    ca_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_227_inst_ack_1, ack => maxPool4_CP_360_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	43 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Sample/rr
      -- CP-element group 136: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Sample/$entry
      -- CP-element group 136: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_sample_start_
      -- 
    rr_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(136), ack => slice_231_inst_req_0); -- 
    maxPool4_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(138);
      gj_maxPool4_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	340 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Update/cr
      -- CP-element group 137: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Update/$entry
      -- CP-element group 137: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_update_start_
      -- 
    cr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(137), ack => slice_231_inst_req_1); -- 
    maxPool4_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(139) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	41 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Sample/ra
      -- CP-element group 138: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_sample_completed_
      -- 
    ra_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_231_inst_ack_0, ack => maxPool4_CP_360_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	338 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Update/ca
      -- CP-element group 139: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_Update/$exit
      -- CP-element group 139: 	 assign_stmt_106_to_assign_stmt_1147/slice_231_update_completed_
      -- 
    ca_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_231_inst_ack_1, ack => maxPool4_CP_360_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	43 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Sample/rr
      -- CP-element group 140: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Sample/$entry
      -- CP-element group 140: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_sample_start_
      -- 
    rr_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(140), ack => slice_235_inst_req_0); -- 
    maxPool4_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(142);
      gj_maxPool4_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	340 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Update/cr
      -- CP-element group 141: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Update/$entry
      -- CP-element group 141: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_update_start_
      -- 
    cr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(141), ack => slice_235_inst_req_1); -- 
    maxPool4_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(143) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	41 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Sample/ra
      -- CP-element group 142: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Sample/$exit
      -- CP-element group 142: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_sample_completed_
      -- 
    ra_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_235_inst_ack_0, ack => maxPool4_CP_360_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	338 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Update/ca
      -- CP-element group 143: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_Update/$exit
      -- CP-element group 143: 	 assign_stmt_106_to_assign_stmt_1147/slice_235_update_completed_
      -- 
    ca_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_235_inst_ack_1, ack => maxPool4_CP_360_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	43 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_sample_start_
      -- CP-element group 144: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Sample/rr
      -- CP-element group 144: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Sample/$entry
      -- 
    rr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(144), ack => slice_239_inst_req_0); -- 
    maxPool4_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(146);
      gj_maxPool4_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	340 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_update_start_
      -- CP-element group 145: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Update/cr
      -- CP-element group 145: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Update/$entry
      -- 
    cr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(145), ack => slice_239_inst_req_1); -- 
    maxPool4_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(147) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	41 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_sample_completed_
      -- CP-element group 146: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Sample/$exit
      -- CP-element group 146: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Sample/ra
      -- 
    ra_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_239_inst_ack_0, ack => maxPool4_CP_360_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	338 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Update/ca
      -- CP-element group 147: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_update_completed_
      -- CP-element group 147: 	 assign_stmt_106_to_assign_stmt_1147/slice_239_Update/$exit
      -- 
    ca_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_239_inst_ack_1, ack => maxPool4_CP_360_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	43 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Sample/rr
      -- CP-element group 148: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Sample/$entry
      -- CP-element group 148: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_sample_start_
      -- 
    rr_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(148), ack => slice_243_inst_req_0); -- 
    maxPool4_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(150);
      gj_maxPool4_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	359 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Update/$entry
      -- CP-element group 149: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_update_start_
      -- CP-element group 149: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Update/cr
      -- 
    cr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(149), ack => slice_243_inst_req_1); -- 
    maxPool4_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(151) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	41 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Sample/ra
      -- CP-element group 150: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Sample/$exit
      -- CP-element group 150: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_sample_completed_
      -- 
    ra_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_243_inst_ack_0, ack => maxPool4_CP_360_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	357 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Update/$exit
      -- CP-element group 151: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_update_completed_
      -- CP-element group 151: 	 assign_stmt_106_to_assign_stmt_1147/slice_243_Update/ca
      -- 
    ca_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_243_inst_ack_1, ack => maxPool4_CP_360_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	43 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Sample/rr
      -- CP-element group 152: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Sample/$entry
      -- CP-element group 152: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_sample_start_
      -- 
    rr_1119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(152), ack => slice_247_inst_req_0); -- 
    maxPool4_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(154);
      gj_maxPool4_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	359 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Update/$entry
      -- CP-element group 153: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_update_start_
      -- CP-element group 153: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Update/cr
      -- 
    cr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(153), ack => slice_247_inst_req_1); -- 
    maxPool4_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(155) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Sample/ra
      -- CP-element group 154: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Sample/$exit
      -- CP-element group 154: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_sample_completed_
      -- 
    ra_1120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_247_inst_ack_0, ack => maxPool4_CP_360_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	357 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Update/$exit
      -- CP-element group 155: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_update_completed_
      -- CP-element group 155: 	 assign_stmt_106_to_assign_stmt_1147/slice_247_Update/ca
      -- 
    ca_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_247_inst_ack_1, ack => maxPool4_CP_360_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	43 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_sample_start_
      -- CP-element group 156: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Sample/rr
      -- CP-element group 156: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Sample/$entry
      -- 
    rr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(156), ack => slice_251_inst_req_0); -- 
    maxPool4_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(158);
      gj_maxPool4_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	359 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Update/$entry
      -- CP-element group 157: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Update/cr
      -- CP-element group 157: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_update_start_
      -- 
    cr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(157), ack => slice_251_inst_req_1); -- 
    maxPool4_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(159) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	41 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Sample/ra
      -- CP-element group 158: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Sample/$exit
      -- CP-element group 158: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_sample_completed_
      -- 
    ra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_251_inst_ack_0, ack => maxPool4_CP_360_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	357 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Update/ca
      -- CP-element group 159: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_update_completed_
      -- CP-element group 159: 	 assign_stmt_106_to_assign_stmt_1147/slice_251_Update/$exit
      -- 
    ca_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_251_inst_ack_1, ack => maxPool4_CP_360_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	43 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Sample/rr
      -- CP-element group 160: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_sample_start_
      -- 
    rr_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(160), ack => slice_255_inst_req_0); -- 
    maxPool4_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(162);
      gj_maxPool4_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	359 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Update/cr
      -- CP-element group 161: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Update/$entry
      -- CP-element group 161: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_update_start_
      -- 
    cr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(161), ack => slice_255_inst_req_1); -- 
    maxPool4_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(163) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	41 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Sample/ra
      -- CP-element group 162: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_sample_completed_
      -- CP-element group 162: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Sample/$exit
      -- 
    ra_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_255_inst_ack_0, ack => maxPool4_CP_360_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	357 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Update/ca
      -- CP-element group 163: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_Update/$exit
      -- CP-element group 163: 	 assign_stmt_106_to_assign_stmt_1147/slice_255_update_completed_
      -- 
    ca_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_255_inst_ack_1, ack => maxPool4_CP_360_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	43 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_sample_start_
      -- CP-element group 164: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Sample/rr
      -- CP-element group 164: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Sample/$entry
      -- 
    rr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(164), ack => slice_259_inst_req_0); -- 
    maxPool4_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(166);
      gj_maxPool4_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	378 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Update/cr
      -- CP-element group 165: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Update/$entry
      -- CP-element group 165: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_update_start_
      -- 
    cr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(165), ack => slice_259_inst_req_1); -- 
    maxPool4_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(167) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	41 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Sample/ra
      -- CP-element group 166: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Sample/$exit
      -- CP-element group 166: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_sample_completed_
      -- 
    ra_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_259_inst_ack_0, ack => maxPool4_CP_360_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	376 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Update/ca
      -- CP-element group 167: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_Update/$exit
      -- CP-element group 167: 	 assign_stmt_106_to_assign_stmt_1147/slice_259_update_completed_
      -- 
    ca_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_259_inst_ack_1, ack => maxPool4_CP_360_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	43 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Sample/$entry
      -- CP-element group 168: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Sample/rr
      -- CP-element group 168: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_sample_start_
      -- 
    rr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(168), ack => slice_263_inst_req_0); -- 
    maxPool4_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(170);
      gj_maxPool4_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	378 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Update/$entry
      -- CP-element group 169: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Update/cr
      -- CP-element group 169: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_update_start_
      -- 
    cr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(169), ack => slice_263_inst_req_1); -- 
    maxPool4_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(171) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	41 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Sample/ra
      -- CP-element group 170: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Sample/$exit
      -- CP-element group 170: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_sample_completed_
      -- 
    ra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_263_inst_ack_0, ack => maxPool4_CP_360_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	376 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Update/ca
      -- CP-element group 171: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_Update/$exit
      -- CP-element group 171: 	 assign_stmt_106_to_assign_stmt_1147/slice_263_update_completed_
      -- 
    ca_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_263_inst_ack_1, ack => maxPool4_CP_360_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	43 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Sample/rr
      -- CP-element group 172: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_sample_start_
      -- 
    rr_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(172), ack => slice_267_inst_req_0); -- 
    maxPool4_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(174);
      gj_maxPool4_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	378 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Update/cr
      -- CP-element group 173: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_update_start_
      -- CP-element group 173: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Update/$entry
      -- 
    cr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(173), ack => slice_267_inst_req_1); -- 
    maxPool4_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(175) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	41 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Sample/$exit
      -- CP-element group 174: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_sample_completed_
      -- CP-element group 174: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Sample/ra
      -- 
    ra_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_267_inst_ack_0, ack => maxPool4_CP_360_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	376 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Update/ca
      -- CP-element group 175: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_update_completed_
      -- CP-element group 175: 	 assign_stmt_106_to_assign_stmt_1147/slice_267_Update/$exit
      -- 
    ca_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_267_inst_ack_1, ack => maxPool4_CP_360_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	43 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_sample_start_
      -- CP-element group 176: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Sample/rr
      -- CP-element group 176: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Sample/$entry
      -- 
    rr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(176), ack => slice_271_inst_req_0); -- 
    maxPool4_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(43) & maxPool4_CP_360_elements(178);
      gj_maxPool4_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	378 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Update/cr
      -- CP-element group 177: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Update/$entry
      -- CP-element group 177: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_update_start_
      -- 
    cr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(177), ack => slice_271_inst_req_1); -- 
    maxPool4_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(179) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	41 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Sample/ra
      -- CP-element group 178: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Sample/$exit
      -- CP-element group 178: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_sample_completed_
      -- 
    ra_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_271_inst_ack_0, ack => maxPool4_CP_360_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	376 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Update/ca
      -- CP-element group 179: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_Update/$exit
      -- CP-element group 179: 	 assign_stmt_106_to_assign_stmt_1147/slice_271_update_completed_
      -- 
    ca_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_271_inst_ack_1, ack => maxPool4_CP_360_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	47 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_sample_start_
      -- CP-element group 180: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Sample/$entry
      -- CP-element group 180: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Sample/rr
      -- 
    rr_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(180), ack => slice_275_inst_req_0); -- 
    maxPool4_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(182);
      gj_maxPool4_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	321 
    -- CP-element group 181: 	386 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Update/cr
      -- CP-element group 181: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Update/$entry
      -- CP-element group 181: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_update_start_
      -- 
    cr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(181), ack => slice_275_inst_req_1); -- 
    maxPool4_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(183) & maxPool4_CP_360_elements(321) & maxPool4_CP_360_elements(386);
      gj_maxPool4_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	45 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_sample_completed_
      -- CP-element group 182: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Sample/$exit
      -- CP-element group 182: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Sample/ra
      -- 
    ra_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_275_inst_ack_0, ack => maxPool4_CP_360_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	319 
    -- CP-element group 183: 	384 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Update/$exit
      -- CP-element group 183: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_update_completed_
      -- CP-element group 183: 	 assign_stmt_106_to_assign_stmt_1147/slice_275_Update/ca
      -- 
    ca_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_275_inst_ack_1, ack => maxPool4_CP_360_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	47 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_sample_start_
      -- CP-element group 184: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Sample/$entry
      -- CP-element group 184: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Sample/rr
      -- 
    rr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(184), ack => slice_279_inst_req_0); -- 
    maxPool4_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(186);
      gj_maxPool4_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	321 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_update_start_
      -- CP-element group 185: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Update/$entry
      -- CP-element group 185: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Update/cr
      -- 
    cr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(185), ack => slice_279_inst_req_1); -- 
    maxPool4_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(187) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	45 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_sample_completed_
      -- CP-element group 186: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Sample/$exit
      -- CP-element group 186: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Sample/ra
      -- 
    ra_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_279_inst_ack_0, ack => maxPool4_CP_360_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	319 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_update_completed_
      -- CP-element group 187: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Update/$exit
      -- CP-element group 187: 	 assign_stmt_106_to_assign_stmt_1147/slice_279_Update/ca
      -- 
    ca_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_279_inst_ack_1, ack => maxPool4_CP_360_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	47 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_sample_start_
      -- CP-element group 188: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Sample/$entry
      -- CP-element group 188: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Sample/rr
      -- 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(188), ack => slice_283_inst_req_0); -- 
    maxPool4_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(190);
      gj_maxPool4_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: 	321 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_update_start_
      -- CP-element group 189: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Update/$entry
      -- CP-element group 189: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Update/cr
      -- 
    cr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(189), ack => slice_283_inst_req_1); -- 
    maxPool4_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(191) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	45 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_sample_completed_
      -- CP-element group 190: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Sample/$exit
      -- CP-element group 190: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Sample/ra
      -- 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_283_inst_ack_0, ack => maxPool4_CP_360_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	319 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_update_completed_
      -- CP-element group 191: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Update/$exit
      -- CP-element group 191: 	 assign_stmt_106_to_assign_stmt_1147/slice_283_Update/ca
      -- 
    ca_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_283_inst_ack_1, ack => maxPool4_CP_360_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	47 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_sample_start_
      -- CP-element group 192: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Sample/$entry
      -- CP-element group 192: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Sample/rr
      -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(192), ack => slice_287_inst_req_0); -- 
    maxPool4_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(194);
      gj_maxPool4_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: 	321 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_update_start_
      -- CP-element group 193: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Update/$entry
      -- CP-element group 193: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Update/cr
      -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(193), ack => slice_287_inst_req_1); -- 
    maxPool4_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(195) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	45 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_sample_completed_
      -- CP-element group 194: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Sample/ra
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_287_inst_ack_0, ack => maxPool4_CP_360_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	319 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_update_completed_
      -- CP-element group 195: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Update/$exit
      -- CP-element group 195: 	 assign_stmt_106_to_assign_stmt_1147/slice_287_Update/ca
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_287_inst_ack_1, ack => maxPool4_CP_360_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	47 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_sample_start_
      -- CP-element group 196: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Sample/$entry
      -- CP-element group 196: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Sample/rr
      -- 
    rr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(196), ack => slice_291_inst_req_0); -- 
    maxPool4_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(198);
      gj_maxPool4_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	340 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_update_start_
      -- CP-element group 197: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Update/$entry
      -- CP-element group 197: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Update/cr
      -- 
    cr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(197), ack => slice_291_inst_req_1); -- 
    maxPool4_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(199) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	45 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_sample_completed_
      -- CP-element group 198: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Sample/$exit
      -- CP-element group 198: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Sample/ra
      -- 
    ra_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_291_inst_ack_0, ack => maxPool4_CP_360_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	338 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_update_completed_
      -- CP-element group 199: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Update/$exit
      -- CP-element group 199: 	 assign_stmt_106_to_assign_stmt_1147/slice_291_Update/ca
      -- 
    ca_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_291_inst_ack_1, ack => maxPool4_CP_360_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	47 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_sample_start_
      -- CP-element group 200: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Sample/$entry
      -- CP-element group 200: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Sample/rr
      -- 
    rr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(200), ack => slice_295_inst_req_0); -- 
    maxPool4_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(202);
      gj_maxPool4_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: 	340 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_update_start_
      -- CP-element group 201: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Update/$entry
      -- CP-element group 201: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Update/cr
      -- 
    cr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(201), ack => slice_295_inst_req_1); -- 
    maxPool4_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(203) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	45 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_sample_completed_
      -- CP-element group 202: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Sample/$exit
      -- CP-element group 202: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Sample/ra
      -- 
    ra_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_295_inst_ack_0, ack => maxPool4_CP_360_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	338 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_update_completed_
      -- CP-element group 203: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Update/$exit
      -- CP-element group 203: 	 assign_stmt_106_to_assign_stmt_1147/slice_295_Update/ca
      -- 
    ca_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_295_inst_ack_1, ack => maxPool4_CP_360_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	47 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_sample_start_
      -- CP-element group 204: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Sample/$entry
      -- CP-element group 204: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Sample/rr
      -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(204), ack => slice_299_inst_req_0); -- 
    maxPool4_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(206);
      gj_maxPool4_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: 	340 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_update_start_
      -- CP-element group 205: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Update/$entry
      -- CP-element group 205: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Update/cr
      -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(205), ack => slice_299_inst_req_1); -- 
    maxPool4_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(207) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	45 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_sample_completed_
      -- CP-element group 206: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Sample/$exit
      -- CP-element group 206: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Sample/ra
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_299_inst_ack_0, ack => maxPool4_CP_360_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	338 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_update_completed_
      -- CP-element group 207: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Update/$exit
      -- CP-element group 207: 	 assign_stmt_106_to_assign_stmt_1147/slice_299_Update/ca
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_299_inst_ack_1, ack => maxPool4_CP_360_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	47 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	210 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_sample_start_
      -- CP-element group 208: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Sample/$entry
      -- CP-element group 208: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Sample/rr
      -- 
    rr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(208), ack => slice_303_inst_req_0); -- 
    maxPool4_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(210);
      gj_maxPool4_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: 	340 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_update_start_
      -- CP-element group 209: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Update/$entry
      -- CP-element group 209: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Update/cr
      -- 
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(209), ack => slice_303_inst_req_1); -- 
    maxPool4_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(211) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_sample_completed_
      -- CP-element group 210: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Sample/$exit
      -- CP-element group 210: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Sample/ra
      -- 
    ra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_303_inst_ack_0, ack => maxPool4_CP_360_elements(210)); -- 
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	338 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_update_completed_
      -- CP-element group 211: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Update/$exit
      -- CP-element group 211: 	 assign_stmt_106_to_assign_stmt_1147/slice_303_Update/ca
      -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_303_inst_ack_1, ack => maxPool4_CP_360_elements(211)); -- 
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	47 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_sample_start_
      -- CP-element group 212: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Sample/$entry
      -- CP-element group 212: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Sample/rr
      -- 
    rr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(212), ack => slice_307_inst_req_0); -- 
    maxPool4_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(214);
      gj_maxPool4_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: 	359 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_update_start_
      -- CP-element group 213: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Update/$entry
      -- CP-element group 213: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Update/cr
      -- 
    cr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(213), ack => slice_307_inst_req_1); -- 
    maxPool4_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(215) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	45 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_sample_completed_
      -- CP-element group 214: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Sample/$exit
      -- CP-element group 214: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Sample/ra
      -- 
    ra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_307_inst_ack_0, ack => maxPool4_CP_360_elements(214)); -- 
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	357 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_update_completed_
      -- CP-element group 215: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Update/$exit
      -- CP-element group 215: 	 assign_stmt_106_to_assign_stmt_1147/slice_307_Update/ca
      -- 
    ca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_307_inst_ack_1, ack => maxPool4_CP_360_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_sample_start_
      -- CP-element group 216: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Sample/$entry
      -- CP-element group 216: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Sample/rr
      -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(216), ack => slice_311_inst_req_0); -- 
    maxPool4_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(218);
      gj_maxPool4_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	359 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_update_start_
      -- CP-element group 217: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Update/$entry
      -- CP-element group 217: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Update/cr
      -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(217), ack => slice_311_inst_req_1); -- 
    maxPool4_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(219) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_sample_completed_
      -- CP-element group 218: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Sample/$exit
      -- CP-element group 218: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Sample/ra
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_311_inst_ack_0, ack => maxPool4_CP_360_elements(218)); -- 
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	357 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_update_completed_
      -- CP-element group 219: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Update/$exit
      -- CP-element group 219: 	 assign_stmt_106_to_assign_stmt_1147/slice_311_Update/ca
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_311_inst_ack_1, ack => maxPool4_CP_360_elements(219)); -- 
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	47 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_sample_start_
      -- CP-element group 220: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Sample/$entry
      -- CP-element group 220: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Sample/rr
      -- 
    rr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(220), ack => slice_315_inst_req_0); -- 
    maxPool4_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(222);
      gj_maxPool4_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: 	359 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_update_start_
      -- CP-element group 221: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Update/$entry
      -- CP-element group 221: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Update/cr
      -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(221), ack => slice_315_inst_req_1); -- 
    maxPool4_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(223) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	45 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_sample_completed_
      -- CP-element group 222: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Sample/$exit
      -- CP-element group 222: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Sample/ra
      -- 
    ra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_315_inst_ack_0, ack => maxPool4_CP_360_elements(222)); -- 
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	357 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_update_completed_
      -- CP-element group 223: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Update/$exit
      -- CP-element group 223: 	 assign_stmt_106_to_assign_stmt_1147/slice_315_Update/ca
      -- 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_315_inst_ack_1, ack => maxPool4_CP_360_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	47 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_sample_start_
      -- CP-element group 224: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Sample/$entry
      -- CP-element group 224: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Sample/rr
      -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(224), ack => slice_319_inst_req_0); -- 
    maxPool4_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(226);
      gj_maxPool4_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: 	359 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_update_start_
      -- CP-element group 225: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Update/$entry
      -- CP-element group 225: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Update/cr
      -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(225), ack => slice_319_inst_req_1); -- 
    maxPool4_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(227) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	45 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_sample_completed_
      -- CP-element group 226: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Sample/$exit
      -- CP-element group 226: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Sample/ra
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_319_inst_ack_0, ack => maxPool4_CP_360_elements(226)); -- 
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	357 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_update_completed_
      -- CP-element group 227: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Update/$exit
      -- CP-element group 227: 	 assign_stmt_106_to_assign_stmt_1147/slice_319_Update/ca
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_319_inst_ack_1, ack => maxPool4_CP_360_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	47 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_sample_start_
      -- CP-element group 228: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Sample/$entry
      -- CP-element group 228: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Sample/rr
      -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(228), ack => slice_323_inst_req_0); -- 
    maxPool4_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(230);
      gj_maxPool4_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	378 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_update_start_
      -- CP-element group 229: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Update/$entry
      -- CP-element group 229: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Update/cr
      -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(229), ack => slice_323_inst_req_1); -- 
    maxPool4_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(231) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	45 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_sample_completed_
      -- CP-element group 230: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Sample/$exit
      -- CP-element group 230: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Sample/ra
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_323_inst_ack_0, ack => maxPool4_CP_360_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	376 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_update_completed_
      -- CP-element group 231: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Update/$exit
      -- CP-element group 231: 	 assign_stmt_106_to_assign_stmt_1147/slice_323_Update/ca
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_323_inst_ack_1, ack => maxPool4_CP_360_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	47 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	234 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_sample_start_
      -- CP-element group 232: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Sample/$entry
      -- CP-element group 232: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Sample/rr
      -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(232), ack => slice_327_inst_req_0); -- 
    maxPool4_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(234);
      gj_maxPool4_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	378 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_update_start_
      -- CP-element group 233: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Update/$entry
      -- CP-element group 233: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Update/cr
      -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(233), ack => slice_327_inst_req_1); -- 
    maxPool4_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(235) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	45 
    -- CP-element group 234: 	232 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_sample_completed_
      -- CP-element group 234: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Sample/$exit
      -- CP-element group 234: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Sample/ra
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_327_inst_ack_0, ack => maxPool4_CP_360_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	376 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_update_completed_
      -- CP-element group 235: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Update/$exit
      -- CP-element group 235: 	 assign_stmt_106_to_assign_stmt_1147/slice_327_Update/ca
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_327_inst_ack_1, ack => maxPool4_CP_360_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	47 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_sample_start_
      -- CP-element group 236: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Sample/$entry
      -- CP-element group 236: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Sample/rr
      -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(236), ack => slice_331_inst_req_0); -- 
    maxPool4_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(238);
      gj_maxPool4_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	378 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_update_start_
      -- CP-element group 237: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Update/$entry
      -- CP-element group 237: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Update/cr
      -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(237), ack => slice_331_inst_req_1); -- 
    maxPool4_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(239) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	45 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_sample_completed_
      -- CP-element group 238: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Sample/$exit
      -- CP-element group 238: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Sample/ra
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_331_inst_ack_0, ack => maxPool4_CP_360_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	376 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_update_completed_
      -- CP-element group 239: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Update/$exit
      -- CP-element group 239: 	 assign_stmt_106_to_assign_stmt_1147/slice_331_Update/ca
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_331_inst_ack_1, ack => maxPool4_CP_360_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	47 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_sample_start_
      -- CP-element group 240: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Sample/$entry
      -- CP-element group 240: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Sample/rr
      -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(240), ack => slice_335_inst_req_0); -- 
    maxPool4_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(47) & maxPool4_CP_360_elements(242);
      gj_maxPool4_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	378 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_update_start_
      -- CP-element group 241: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Update/$entry
      -- CP-element group 241: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Update/cr
      -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(241), ack => slice_335_inst_req_1); -- 
    maxPool4_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(243) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	45 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_sample_completed_
      -- CP-element group 242: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Sample/$exit
      -- CP-element group 242: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Sample/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_335_inst_ack_0, ack => maxPool4_CP_360_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	376 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_update_completed_
      -- CP-element group 243: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Update/$exit
      -- CP-element group 243: 	 assign_stmt_106_to_assign_stmt_1147/slice_335_Update/ca
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_335_inst_ack_1, ack => maxPool4_CP_360_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	51 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_sample_start_
      -- CP-element group 244: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Sample/$entry
      -- CP-element group 244: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Sample/rr
      -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(244), ack => slice_339_inst_req_0); -- 
    maxPool4_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(246);
      gj_maxPool4_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	321 
    -- CP-element group 245: 	386 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_update_start_
      -- CP-element group 245: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Update/$entry
      -- CP-element group 245: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Update/cr
      -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(245), ack => slice_339_inst_req_1); -- 
    maxPool4_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(247) & maxPool4_CP_360_elements(321) & maxPool4_CP_360_elements(386);
      gj_maxPool4_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	49 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_sample_completed_
      -- CP-element group 246: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Sample/$exit
      -- CP-element group 246: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Sample/ra
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_339_inst_ack_0, ack => maxPool4_CP_360_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	319 
    -- CP-element group 247: 	384 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_update_completed_
      -- CP-element group 247: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Update/$exit
      -- CP-element group 247: 	 assign_stmt_106_to_assign_stmt_1147/slice_339_Update/ca
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_339_inst_ack_1, ack => maxPool4_CP_360_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	51 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_sample_start_
      -- CP-element group 248: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Sample/$entry
      -- CP-element group 248: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Sample/rr
      -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(248), ack => slice_343_inst_req_0); -- 
    maxPool4_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(250);
      gj_maxPool4_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	321 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_update_start_
      -- CP-element group 249: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Update/$entry
      -- CP-element group 249: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Update/cr
      -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(249), ack => slice_343_inst_req_1); -- 
    maxPool4_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(251) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	49 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_sample_completed_
      -- CP-element group 250: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Sample/$exit
      -- CP-element group 250: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Sample/ra
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_343_inst_ack_0, ack => maxPool4_CP_360_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	319 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_update_completed_
      -- CP-element group 251: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Update/$exit
      -- CP-element group 251: 	 assign_stmt_106_to_assign_stmt_1147/slice_343_Update/ca
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_343_inst_ack_1, ack => maxPool4_CP_360_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	51 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_sample_start_
      -- CP-element group 252: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Sample/$entry
      -- CP-element group 252: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Sample/rr
      -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(252), ack => slice_347_inst_req_0); -- 
    maxPool4_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(254);
      gj_maxPool4_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	321 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_update_start_
      -- CP-element group 253: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Update/$entry
      -- CP-element group 253: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Update/cr
      -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(253), ack => slice_347_inst_req_1); -- 
    maxPool4_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(255) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	49 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_sample_completed_
      -- CP-element group 254: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Sample/$exit
      -- CP-element group 254: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Sample/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_347_inst_ack_0, ack => maxPool4_CP_360_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	319 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_update_completed_
      -- CP-element group 255: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Update/$exit
      -- CP-element group 255: 	 assign_stmt_106_to_assign_stmt_1147/slice_347_Update/ca
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_347_inst_ack_1, ack => maxPool4_CP_360_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	51 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_sample_start_
      -- CP-element group 256: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Sample/$entry
      -- CP-element group 256: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Sample/rr
      -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(256), ack => slice_351_inst_req_0); -- 
    maxPool4_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(258);
      gj_maxPool4_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	321 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_update_start_
      -- CP-element group 257: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Update/$entry
      -- CP-element group 257: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Update/cr
      -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(257), ack => slice_351_inst_req_1); -- 
    maxPool4_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(259) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	49 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_sample_completed_
      -- CP-element group 258: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Sample/$exit
      -- CP-element group 258: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Sample/ra
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_351_inst_ack_0, ack => maxPool4_CP_360_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	319 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_update_completed_
      -- CP-element group 259: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Update/$exit
      -- CP-element group 259: 	 assign_stmt_106_to_assign_stmt_1147/slice_351_Update/ca
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_351_inst_ack_1, ack => maxPool4_CP_360_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	51 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_sample_start_
      -- CP-element group 260: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Sample/$entry
      -- CP-element group 260: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Sample/rr
      -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(260), ack => slice_355_inst_req_0); -- 
    maxPool4_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(262);
      gj_maxPool4_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	340 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_update_start_
      -- CP-element group 261: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Update/$entry
      -- CP-element group 261: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Update/cr
      -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(261), ack => slice_355_inst_req_1); -- 
    maxPool4_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(263) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	49 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_sample_completed_
      -- CP-element group 262: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Sample/$exit
      -- CP-element group 262: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_355_inst_ack_0, ack => maxPool4_CP_360_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	338 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_update_completed_
      -- CP-element group 263: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Update/$exit
      -- CP-element group 263: 	 assign_stmt_106_to_assign_stmt_1147/slice_355_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_355_inst_ack_1, ack => maxPool4_CP_360_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	51 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_sample_start_
      -- CP-element group 264: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Sample/$entry
      -- CP-element group 264: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Sample/rr
      -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(264), ack => slice_359_inst_req_0); -- 
    maxPool4_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(266);
      gj_maxPool4_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: 	340 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_update_start_
      -- CP-element group 265: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Update/$entry
      -- CP-element group 265: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Update/cr
      -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(265), ack => slice_359_inst_req_1); -- 
    maxPool4_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(267) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	49 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_sample_completed_
      -- CP-element group 266: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Sample/$exit
      -- CP-element group 266: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Sample/ra
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_359_inst_ack_0, ack => maxPool4_CP_360_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	338 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_update_completed_
      -- CP-element group 267: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Update/$exit
      -- CP-element group 267: 	 assign_stmt_106_to_assign_stmt_1147/slice_359_Update/ca
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_359_inst_ack_1, ack => maxPool4_CP_360_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	51 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_sample_start_
      -- CP-element group 268: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Sample/$entry
      -- CP-element group 268: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Sample/rr
      -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(268), ack => slice_363_inst_req_0); -- 
    maxPool4_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(270);
      gj_maxPool4_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	340 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_update_start_
      -- CP-element group 269: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Update/$entry
      -- CP-element group 269: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Update/cr
      -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(269), ack => slice_363_inst_req_1); -- 
    maxPool4_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(271) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	49 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_sample_completed_
      -- CP-element group 270: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Sample/$exit
      -- CP-element group 270: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Sample/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_363_inst_ack_0, ack => maxPool4_CP_360_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	338 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_update_completed_
      -- CP-element group 271: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Update/$exit
      -- CP-element group 271: 	 assign_stmt_106_to_assign_stmt_1147/slice_363_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_363_inst_ack_1, ack => maxPool4_CP_360_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	51 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_sample_start_
      -- CP-element group 272: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Sample/$entry
      -- CP-element group 272: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Sample/rr
      -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(272), ack => slice_367_inst_req_0); -- 
    maxPool4_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(274);
      gj_maxPool4_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	340 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_update_start_
      -- CP-element group 273: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Update/$entry
      -- CP-element group 273: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Update/cr
      -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(273), ack => slice_367_inst_req_1); -- 
    maxPool4_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(275) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	49 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_sample_completed_
      -- CP-element group 274: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Sample/$exit
      -- CP-element group 274: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Sample/ra
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_367_inst_ack_0, ack => maxPool4_CP_360_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	338 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_update_completed_
      -- CP-element group 275: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Update/$exit
      -- CP-element group 275: 	 assign_stmt_106_to_assign_stmt_1147/slice_367_Update/ca
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_367_inst_ack_1, ack => maxPool4_CP_360_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	51 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_sample_start_
      -- CP-element group 276: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Sample/$entry
      -- CP-element group 276: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Sample/rr
      -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(276), ack => slice_371_inst_req_0); -- 
    maxPool4_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(278);
      gj_maxPool4_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: 	359 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_update_start_
      -- CP-element group 277: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Update/$entry
      -- CP-element group 277: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Update/cr
      -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(277), ack => slice_371_inst_req_1); -- 
    maxPool4_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(279) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	49 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_sample_completed_
      -- CP-element group 278: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Sample/$exit
      -- CP-element group 278: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Sample/ra
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_371_inst_ack_0, ack => maxPool4_CP_360_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	357 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_update_completed_
      -- CP-element group 279: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Update/$exit
      -- CP-element group 279: 	 assign_stmt_106_to_assign_stmt_1147/slice_371_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_371_inst_ack_1, ack => maxPool4_CP_360_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	51 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Sample/rr
      -- CP-element group 280: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Sample/$entry
      -- CP-element group 280: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_sample_start_
      -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(280), ack => slice_375_inst_req_0); -- 
    maxPool4_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(282);
      gj_maxPool4_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: 	359 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Update/cr
      -- CP-element group 281: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Update/$entry
      -- CP-element group 281: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_update_start_
      -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(281), ack => slice_375_inst_req_1); -- 
    maxPool4_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(283) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	49 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Sample/ra
      -- CP-element group 282: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Sample/$exit
      -- CP-element group 282: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_sample_completed_
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_375_inst_ack_0, ack => maxPool4_CP_360_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	357 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Update/ca
      -- CP-element group 283: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_Update/$exit
      -- CP-element group 283: 	 assign_stmt_106_to_assign_stmt_1147/slice_375_update_completed_
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_375_inst_ack_1, ack => maxPool4_CP_360_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	51 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Sample/rr
      -- CP-element group 284: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Sample/$entry
      -- CP-element group 284: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_sample_start_
      -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(284), ack => slice_379_inst_req_0); -- 
    maxPool4_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(286);
      gj_maxPool4_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	359 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Update/cr
      -- CP-element group 285: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Update/$entry
      -- CP-element group 285: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_update_start_
      -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(285), ack => slice_379_inst_req_1); -- 
    maxPool4_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(287) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	49 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Sample/$exit
      -- CP-element group 286: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Sample/ra
      -- CP-element group 286: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_sample_completed_
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_379_inst_ack_0, ack => maxPool4_CP_360_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	357 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Update/$exit
      -- CP-element group 287: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_Update/ca
      -- CP-element group 287: 	 assign_stmt_106_to_assign_stmt_1147/slice_379_update_completed_
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_379_inst_ack_1, ack => maxPool4_CP_360_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	51 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_sample_start_
      -- CP-element group 288: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Sample/rr
      -- CP-element group 288: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Sample/$entry
      -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(288), ack => slice_383_inst_req_0); -- 
    maxPool4_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(290);
      gj_maxPool4_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: 	359 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_update_start_
      -- CP-element group 289: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Update/$entry
      -- CP-element group 289: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Update/cr
      -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(289), ack => slice_383_inst_req_1); -- 
    maxPool4_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(291) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	49 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_sample_completed_
      -- CP-element group 290: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Sample/ra
      -- CP-element group 290: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Sample/$exit
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_383_inst_ack_0, ack => maxPool4_CP_360_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	357 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_update_completed_
      -- CP-element group 291: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Update/$exit
      -- CP-element group 291: 	 assign_stmt_106_to_assign_stmt_1147/slice_383_Update/ca
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_383_inst_ack_1, ack => maxPool4_CP_360_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	51 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Sample/rr
      -- CP-element group 292: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Sample/$entry
      -- CP-element group 292: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_sample_start_
      -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(292), ack => slice_387_inst_req_0); -- 
    maxPool4_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(294);
      gj_maxPool4_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: 	378 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Update/$entry
      -- CP-element group 293: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Update/cr
      -- CP-element group 293: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_update_start_
      -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(293), ack => slice_387_inst_req_1); -- 
    maxPool4_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(295) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	49 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Sample/$exit
      -- CP-element group 294: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Sample/ra
      -- CP-element group 294: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_sample_completed_
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_387_inst_ack_0, ack => maxPool4_CP_360_elements(294)); -- 
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	376 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_update_completed_
      -- CP-element group 295: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Update/$exit
      -- CP-element group 295: 	 assign_stmt_106_to_assign_stmt_1147/slice_387_Update/ca
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_387_inst_ack_1, ack => maxPool4_CP_360_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	51 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	298 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_sample_start_
      -- CP-element group 296: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Sample/rr
      -- CP-element group 296: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Sample/$entry
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(296), ack => slice_391_inst_req_0); -- 
    maxPool4_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(298);
      gj_maxPool4_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: 	378 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_update_start_
      -- CP-element group 297: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Update/cr
      -- CP-element group 297: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Update/$entry
      -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(297), ack => slice_391_inst_req_1); -- 
    maxPool4_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(299) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: marked-successors 
    -- CP-element group 298: 	49 
    -- CP-element group 298: 	296 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_sample_completed_
      -- CP-element group 298: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Sample/ra
      -- CP-element group 298: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Sample/$exit
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_391_inst_ack_0, ack => maxPool4_CP_360_elements(298)); -- 
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	376 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_update_completed_
      -- CP-element group 299: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Update/ca
      -- CP-element group 299: 	 assign_stmt_106_to_assign_stmt_1147/slice_391_Update/$exit
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_391_inst_ack_1, ack => maxPool4_CP_360_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	51 
    -- CP-element group 300: marked-predecessors 
    -- CP-element group 300: 	302 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Sample/rr
      -- CP-element group 300: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Sample/$entry
      -- CP-element group 300: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_sample_start_
      -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(300), ack => slice_395_inst_req_0); -- 
    maxPool4_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(302);
      gj_maxPool4_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: 	378 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Update/cr
      -- CP-element group 301: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Update/$entry
      -- CP-element group 301: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_update_start_
      -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(301), ack => slice_395_inst_req_1); -- 
    maxPool4_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(303) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: successors 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	49 
    -- CP-element group 302: 	300 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Sample/ra
      -- CP-element group 302: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Sample/$exit
      -- CP-element group 302: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_sample_completed_
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_395_inst_ack_0, ack => maxPool4_CP_360_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	376 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Update/ca
      -- CP-element group 303: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_Update/$exit
      -- CP-element group 303: 	 assign_stmt_106_to_assign_stmt_1147/slice_395_update_completed_
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_395_inst_ack_1, ack => maxPool4_CP_360_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	51 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Sample/$entry
      -- CP-element group 304: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_sample_start_
      -- CP-element group 304: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Sample/rr
      -- 
    rr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(304), ack => slice_399_inst_req_0); -- 
    maxPool4_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(51) & maxPool4_CP_360_elements(306);
      gj_maxPool4_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	378 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Update/$entry
      -- CP-element group 305: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_update_start_
      -- CP-element group 305: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Update/cr
      -- 
    cr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(305), ack => slice_399_inst_req_1); -- 
    maxPool4_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(307) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: marked-successors 
    -- CP-element group 306: 	49 
    -- CP-element group 306: 	304 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Sample/ra
      -- CP-element group 306: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_sample_completed_
      -- CP-element group 306: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Sample/$exit
      -- 
    ra_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_399_inst_ack_0, ack => maxPool4_CP_360_elements(306)); -- 
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	376 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Update/$exit
      -- CP-element group 307: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_Update/ca
      -- CP-element group 307: 	 assign_stmt_106_to_assign_stmt_1147/slice_399_update_completed_
      -- 
    ca_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_399_inst_ack_1, ack => maxPool4_CP_360_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	312 
    -- CP-element group 308: marked-predecessors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_request/$entry
      -- CP-element group 308: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_request/req
      -- CP-element group 308: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_sample_start_
      -- 
    req_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(308), ack => addr_of_1047_final_reg_req_0); -- 
    maxPool4_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(312) & maxPool4_CP_360_elements(313);
      gj_maxPool4_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	1 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: 	317 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	314 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_complete/$entry
      -- CP-element group 309: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_update_start_
      -- CP-element group 309: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_complete/req
      -- 
    req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(309), ack => addr_of_1047_final_reg_req_1); -- 
    maxPool4_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(314) & maxPool4_CP_360_elements(317);
      gj_maxPool4_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	1 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	313 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_update_start
      -- CP-element group 310: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Update/$entry
      -- CP-element group 310: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Update/req
      -- 
    req_1687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(310), ack => array_obj_ref_1046_index_offset_req_1); -- 
    maxPool4_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(312) & maxPool4_CP_360_elements(313);
      gj_maxPool4_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	1 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	391 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	2 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_sample_complete
      -- CP-element group 311: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Sample/$exit
      -- CP-element group 311: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Sample/ack
      -- 
    ack_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_offset_ack_0, ack => maxPool4_CP_360_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (8) 
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_base_plus_offset/sum_rename_req
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_base_plus_offset/sum_rename_ack
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_base_plus_offset/$entry
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_base_plus_offset/$exit
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_root_address_calculated
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_offset_calculated
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Update/$exit
      -- CP-element group 312: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1046_final_index_sum_regn_Update/ack
      -- 
    ack_1688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1046_index_offset_ack_1, ack => maxPool4_CP_360_elements(312)); -- 
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: successors 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	310 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_request/ack
      -- CP-element group 313: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_request/$exit
      -- CP-element group 313: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_sample_completed_
      -- 
    ack_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1047_final_reg_ack_0, ack => maxPool4_CP_360_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_complete/$exit
      -- CP-element group 314: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_update_completed_
      -- CP-element group 314: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1047_complete/ack
      -- 
    ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1047_final_reg_ack_1, ack => maxPool4_CP_360_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_sample_start_
      -- CP-element group 315: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Sample/$entry
      -- CP-element group 315: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Sample/req
      -- 
    req_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(315), ack => W_myptr5_1049_delayed_8_0_1049_inst_req_0); -- 
    maxPool4_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(314) & maxPool4_CP_360_elements(317);
      gj_maxPool4_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: marked-predecessors 
    -- CP-element group 316: 	318 
    -- CP-element group 316: 	325 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Update/$entry
      -- CP-element group 316: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Update/req
      -- CP-element group 316: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_update_start_
      -- 
    req_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(316), ack => W_myptr5_1049_delayed_8_0_1049_inst_req_1); -- 
    maxPool4_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(318) & maxPool4_CP_360_elements(325);
      gj_maxPool4_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: marked-successors 
    -- CP-element group 317: 	309 
    -- CP-element group 317: 	315 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Sample/ack
      -- CP-element group 317: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_sample_completed_
      -- CP-element group 317: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Sample/$exit
      -- 
    ack_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1049_delayed_8_0_1049_inst_ack_0, ack => maxPool4_CP_360_elements(317)); -- 
    -- CP-element group 318:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	323 
    -- CP-element group 318: marked-successors 
    -- CP-element group 318: 	316 
    -- CP-element group 318:  members (19) 
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Update/ack
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_Update/$exit
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_address_calculated
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_word_address_calculated
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_root_address_calculated
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_address_resized
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_addr_resize/$entry
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_addr_resize/$exit
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_addr_resize/base_resize_req
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_addr_resize/base_resize_ack
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_plus_offset/$entry
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_plus_offset/$exit
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_plus_offset/sum_rename_req
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_base_plus_offset/sum_rename_ack
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_word_addrgen/$entry
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_word_addrgen/$exit
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_word_addrgen/root_register_req
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_word_addrgen/root_register_ack
      -- CP-element group 318: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1051_update_completed_
      -- 
    ack_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1049_delayed_8_0_1049_inst_ack_1, ack => maxPool4_CP_360_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	55 
    -- CP-element group 319: 	59 
    -- CP-element group 319: 	63 
    -- CP-element group 319: 	67 
    -- CP-element group 319: 	119 
    -- CP-element group 319: 	123 
    -- CP-element group 319: 	127 
    -- CP-element group 319: 	131 
    -- CP-element group 319: 	183 
    -- CP-element group 319: 	187 
    -- CP-element group 319: 	191 
    -- CP-element group 319: 	195 
    -- CP-element group 319: 	247 
    -- CP-element group 319: 	251 
    -- CP-element group 319: 	255 
    -- CP-element group 319: 	259 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Sample/$entry
      -- CP-element group 319: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_sample_start_
      -- CP-element group 319: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Sample/rr
      -- 
    rr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(319), ack => CONCAT_u32_u64_1064_inst_req_0); -- 
    maxPool4_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(55) & maxPool4_CP_360_elements(59) & maxPool4_CP_360_elements(63) & maxPool4_CP_360_elements(67) & maxPool4_CP_360_elements(119) & maxPool4_CP_360_elements(123) & maxPool4_CP_360_elements(127) & maxPool4_CP_360_elements(131) & maxPool4_CP_360_elements(183) & maxPool4_CP_360_elements(187) & maxPool4_CP_360_elements(191) & maxPool4_CP_360_elements(195) & maxPool4_CP_360_elements(247) & maxPool4_CP_360_elements(251) & maxPool4_CP_360_elements(255) & maxPool4_CP_360_elements(259) & maxPool4_CP_360_elements(321);
      gj_maxPool4_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: marked-predecessors 
    -- CP-element group 320: 	322 
    -- CP-element group 320: 	325 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_update_start_
      -- CP-element group 320: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Update/$entry
      -- CP-element group 320: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Update/cr
      -- 
    cr_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(320), ack => CONCAT_u32_u64_1064_inst_req_1); -- 
    maxPool4_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(322) & maxPool4_CP_360_elements(325);
      gj_maxPool4_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	53 
    -- CP-element group 321: 	57 
    -- CP-element group 321: 	61 
    -- CP-element group 321: 	65 
    -- CP-element group 321: 	117 
    -- CP-element group 321: 	121 
    -- CP-element group 321: 	125 
    -- CP-element group 321: 	129 
    -- CP-element group 321: 	181 
    -- CP-element group 321: 	185 
    -- CP-element group 321: 	189 
    -- CP-element group 321: 	193 
    -- CP-element group 321: 	245 
    -- CP-element group 321: 	249 
    -- CP-element group 321: 	253 
    -- CP-element group 321: 	257 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Sample/ra
      -- CP-element group 321: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Sample/$exit
      -- CP-element group 321: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_sample_completed_
      -- 
    ra_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1064_inst_ack_0, ack => maxPool4_CP_360_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322: marked-successors 
    -- CP-element group 322: 	320 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_update_completed_
      -- CP-element group 322: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Update/$exit
      -- CP-element group 322: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1064_Update/ca
      -- 
    ca_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1064_inst_ack_1, ack => maxPool4_CP_360_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	322 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	325 
    -- CP-element group 323: 	382 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (9) 
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_sample_start_
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/$entry
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/ptr_deref_1053_Split/$entry
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/ptr_deref_1053_Split/$exit
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/ptr_deref_1053_Split/split_req
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/ptr_deref_1053_Split/split_ack
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/$entry
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/word_0/$entry
      -- CP-element group 323: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/word_0/rr
      -- 
    rr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(323), ack => ptr_deref_1053_store_0_req_0); -- 
    maxPool4_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(318) & maxPool4_CP_360_elements(322) & maxPool4_CP_360_elements(325) & maxPool4_CP_360_elements(382);
      gj_maxPool4_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: marked-predecessors 
    -- CP-element group 324: 	326 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/$entry
      -- CP-element group 324: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/word_0/cr
      -- CP-element group 324: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/word_0/$entry
      -- CP-element group 324: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_update_start_
      -- CP-element group 324: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/$entry
      -- 
    cr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(324), ack => ptr_deref_1053_store_0_req_1); -- 
    maxPool4_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(326);
      gj_maxPool4_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	388 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	316 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	323 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/$exit
      -- CP-element group 325: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_sample_completed_
      -- CP-element group 325: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/$exit
      -- CP-element group 325: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/word_0/$exit
      -- CP-element group 325: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Sample/word_access_start/word_0/ra
      -- 
    ra_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1053_store_0_ack_0, ack => maxPool4_CP_360_elements(325)); -- 
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	391 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	324 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/$exit
      -- CP-element group 326: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/word_0/ca
      -- CP-element group 326: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/word_access_complete/word_0/$exit
      -- CP-element group 326: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_update_completed_
      -- CP-element group 326: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_Update/$exit
      -- 
    ca_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1053_store_0_ack_1, ack => maxPool4_CP_360_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	331 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	332 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	332 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_request/$entry
      -- CP-element group 327: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_sample_start_
      -- CP-element group 327: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_request/req
      -- 
    req_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(327), ack => addr_of_1073_final_reg_req_0); -- 
    maxPool4_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(331) & maxPool4_CP_360_elements(332);
      gj_maxPool4_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	1 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	333 
    -- CP-element group 328: 	336 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	333 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_update_start_
      -- CP-element group 328: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_complete/$entry
      -- CP-element group 328: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_complete/req
      -- 
    req_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(328), ack => addr_of_1073_final_reg_req_1); -- 
    maxPool4_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(333) & maxPool4_CP_360_elements(336);
      gj_maxPool4_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	1 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: 	332 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Update/$entry
      -- CP-element group 329: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Update/req
      -- CP-element group 329: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_update_start
      -- 
    req_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(329), ack => array_obj_ref_1072_index_offset_req_1); -- 
    maxPool4_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(331) & maxPool4_CP_360_elements(332);
      gj_maxPool4_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	1 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	391 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	2 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_sample_complete
      -- CP-element group 330: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Sample/$exit
      -- CP-element group 330: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Sample/ack
      -- 
    ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_0, ack => maxPool4_CP_360_elements(330)); -- 
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	327 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (8) 
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Update/$exit
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_final_index_sum_regn_Update/ack
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_root_address_calculated
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_offset_calculated
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_base_plus_offset/$entry
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_base_plus_offset/sum_rename_req
      -- CP-element group 331: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1072_base_plus_offset/$exit
      -- 
    ack_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1072_index_offset_ack_1, ack => maxPool4_CP_360_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: 	329 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_sample_completed_
      -- CP-element group 332: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_request/$exit
      -- CP-element group 332: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_request/ack
      -- 
    ack_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_0, ack => maxPool4_CP_360_elements(332)); -- 
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	328 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	328 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_complete/ack
      -- CP-element group 333: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_update_completed_
      -- CP-element group 333: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1073_complete/$exit
      -- 
    ack_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1073_final_reg_ack_1, ack => maxPool4_CP_360_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Sample/req
      -- CP-element group 334: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Sample/$entry
      -- CP-element group 334: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_sample_start_
      -- 
    req_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(334), ack => W_myptr6_1072_delayed_8_0_1075_inst_req_0); -- 
    maxPool4_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(333) & maxPool4_CP_360_elements(336);
      gj_maxPool4_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	344 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Update/$entry
      -- CP-element group 335: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Update/req
      -- CP-element group 335: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_update_start_
      -- 
    req_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(335), ack => W_myptr6_1072_delayed_8_0_1075_inst_req_1); -- 
    maxPool4_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(337) & maxPool4_CP_360_elements(344);
      gj_maxPool4_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Sample/ack
      -- CP-element group 336: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Sample/$exit
      -- CP-element group 336: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_sample_completed_
      -- 
    ack_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1072_delayed_8_0_1075_inst_ack_0, ack => maxPool4_CP_360_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Update/$exit
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_addr_resize/$entry
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_addr_resize/$exit
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_address_calculated
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_plus_offset/sum_rename_req
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_word_addrgen/$entry
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_word_addrgen/$exit
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_plus_offset/$entry
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_plus_offset/$exit
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_Update/ack
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_root_address_calculated
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_address_resized
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_word_address_calculated
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_word_addrgen/root_register_ack
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_word_addrgen/root_register_req
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1077_update_completed_
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_base_addr_resize/base_resize_req
      -- 
    ack_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1072_delayed_8_0_1075_inst_ack_1, ack => maxPool4_CP_360_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	71 
    -- CP-element group 338: 	75 
    -- CP-element group 338: 	79 
    -- CP-element group 338: 	83 
    -- CP-element group 338: 	135 
    -- CP-element group 338: 	139 
    -- CP-element group 338: 	143 
    -- CP-element group 338: 	147 
    -- CP-element group 338: 	199 
    -- CP-element group 338: 	203 
    -- CP-element group 338: 	207 
    -- CP-element group 338: 	211 
    -- CP-element group 338: 	263 
    -- CP-element group 338: 	267 
    -- CP-element group 338: 	271 
    -- CP-element group 338: 	275 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Sample/rr
      -- CP-element group 338: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Sample/$entry
      -- CP-element group 338: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_sample_start_
      -- 
    rr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(338), ack => CONCAT_u32_u64_1090_inst_req_0); -- 
    maxPool4_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(71) & maxPool4_CP_360_elements(75) & maxPool4_CP_360_elements(79) & maxPool4_CP_360_elements(83) & maxPool4_CP_360_elements(135) & maxPool4_CP_360_elements(139) & maxPool4_CP_360_elements(143) & maxPool4_CP_360_elements(147) & maxPool4_CP_360_elements(199) & maxPool4_CP_360_elements(203) & maxPool4_CP_360_elements(207) & maxPool4_CP_360_elements(211) & maxPool4_CP_360_elements(263) & maxPool4_CP_360_elements(267) & maxPool4_CP_360_elements(271) & maxPool4_CP_360_elements(275) & maxPool4_CP_360_elements(340);
      gj_maxPool4_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	344 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Update/$entry
      -- CP-element group 339: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_update_start_
      -- CP-element group 339: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Update/cr
      -- 
    cr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(339), ack => CONCAT_u32_u64_1090_inst_req_1); -- 
    maxPool4_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(341) & maxPool4_CP_360_elements(344);
      gj_maxPool4_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	69 
    -- CP-element group 340: 	73 
    -- CP-element group 340: 	77 
    -- CP-element group 340: 	81 
    -- CP-element group 340: 	133 
    -- CP-element group 340: 	137 
    -- CP-element group 340: 	141 
    -- CP-element group 340: 	145 
    -- CP-element group 340: 	197 
    -- CP-element group 340: 	201 
    -- CP-element group 340: 	205 
    -- CP-element group 340: 	209 
    -- CP-element group 340: 	261 
    -- CP-element group 340: 	265 
    -- CP-element group 340: 	269 
    -- CP-element group 340: 	273 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Sample/$exit
      -- CP-element group 340: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Sample/ra
      -- CP-element group 340: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_sample_completed_
      -- 
    ra_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1090_inst_ack_0, ack => maxPool4_CP_360_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Update/$exit
      -- CP-element group 341: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_update_completed_
      -- CP-element group 341: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1090_Update/ca
      -- 
    ca_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1090_inst_ack_1, ack => maxPool4_CP_360_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: 	341 
    -- CP-element group 342: 	388 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (9) 
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/ptr_deref_1079_Split/$exit
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/ptr_deref_1079_Split/split_req
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/ptr_deref_1079_Split/split_ack
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/$entry
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_sample_start_
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/ptr_deref_1079_Split/$entry
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/$entry
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/word_0/$entry
      -- CP-element group 342: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/word_0/rr
      -- 
    rr_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(342), ack => ptr_deref_1079_store_0_req_0); -- 
    maxPool4_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(337) & maxPool4_CP_360_elements(341) & maxPool4_CP_360_elements(388) & maxPool4_CP_360_elements(344);
      gj_maxPool4_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_update_start_
      -- CP-element group 343: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/$entry
      -- CP-element group 343: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/$entry
      -- CP-element group 343: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/word_0/cr
      -- 
    cr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(343), ack => ptr_deref_1079_store_0_req_1); -- 
    maxPool4_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(345);
      gj_maxPool4_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	389 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: 	339 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_sample_completed_
      -- CP-element group 344: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/$exit
      -- CP-element group 344: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/$exit
      -- CP-element group 344: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/word_0/$exit
      -- CP-element group 344: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Sample/word_access_start/word_0/ra
      -- 
    ra_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1079_store_0_ack_0, ack => maxPool4_CP_360_elements(344)); -- 
    -- CP-element group 345:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	391 
    -- CP-element group 345: marked-successors 
    -- CP-element group 345: 	343 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_update_completed_
      -- CP-element group 345: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/$exit
      -- CP-element group 345: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/$exit
      -- CP-element group 345: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/word_0/$exit
      -- CP-element group 345: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_Update/word_access_complete/word_0/ca
      -- 
    ca_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1079_store_0_ack_1, ack => maxPool4_CP_360_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	350 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	351 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_sample_start_
      -- CP-element group 346: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_request/$entry
      -- CP-element group 346: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_request/req
      -- 
    req_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(346), ack => addr_of_1099_final_reg_req_0); -- 
    maxPool4_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(350) & maxPool4_CP_360_elements(351);
      gj_maxPool4_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	1 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	352 
    -- CP-element group 347: 	355 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	352 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_update_start_
      -- CP-element group 347: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_complete/$entry
      -- CP-element group 347: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_complete/req
      -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(347), ack => addr_of_1099_final_reg_req_1); -- 
    maxPool4_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(352) & maxPool4_CP_360_elements(355);
      gj_maxPool4_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	1 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	351 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_update_start
      -- CP-element group 348: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Update/$entry
      -- CP-element group 348: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Update/req
      -- 
    req_1935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(348), ack => array_obj_ref_1098_index_offset_req_1); -- 
    maxPool4_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(350) & maxPool4_CP_360_elements(351);
      gj_maxPool4_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	1 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	391 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	2 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_sample_complete
      -- CP-element group 349: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Sample/$exit
      -- CP-element group 349: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Sample/ack
      -- 
    ack_1931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_index_offset_ack_0, ack => maxPool4_CP_360_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	346 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (8) 
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_root_address_calculated
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_offset_calculated
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Update/$exit
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_final_index_sum_regn_Update/ack
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_base_plus_offset/$entry
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_base_plus_offset/$exit
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_base_plus_offset/sum_rename_req
      -- CP-element group 350: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1098_base_plus_offset/sum_rename_ack
      -- 
    ack_1936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1098_index_offset_ack_1, ack => maxPool4_CP_360_elements(350)); -- 
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	348 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_sample_completed_
      -- CP-element group 351: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_request/$exit
      -- CP-element group 351: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_request/ack
      -- 
    ack_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1099_final_reg_ack_0, ack => maxPool4_CP_360_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	347 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	347 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_update_completed_
      -- CP-element group 352: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_complete/$exit
      -- CP-element group 352: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1099_complete/ack
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1099_final_reg_ack_1, ack => maxPool4_CP_360_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_sample_start_
      -- CP-element group 353: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Sample/$entry
      -- CP-element group 353: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Sample/req
      -- 
    req_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(353), ack => W_myptr7_1095_delayed_8_0_1101_inst_req_0); -- 
    maxPool4_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(352) & maxPool4_CP_360_elements(355);
      gj_maxPool4_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: 	363 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_update_start_
      -- CP-element group 354: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Update/$entry
      -- CP-element group 354: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Update/req
      -- 
    req_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(354), ack => W_myptr7_1095_delayed_8_0_1101_inst_req_1); -- 
    maxPool4_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(356) & maxPool4_CP_360_elements(363);
      gj_maxPool4_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	347 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_sample_completed_
      -- CP-element group 355: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Sample/$exit
      -- CP-element group 355: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Sample/ack
      -- 
    ack_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1095_delayed_8_0_1101_inst_ack_0, ack => maxPool4_CP_360_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	361 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (19) 
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_update_completed_
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Update/$exit
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1103_Update/ack
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_address_calculated
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_word_address_calculated
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_root_address_calculated
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_address_resized
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_addr_resize/$entry
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_addr_resize/$exit
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_addr_resize/base_resize_req
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_addr_resize/base_resize_ack
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_plus_offset/$entry
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_plus_offset/$exit
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_plus_offset/sum_rename_req
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_base_plus_offset/sum_rename_ack
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_word_addrgen/$entry
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_word_addrgen/$exit
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_word_addrgen/root_register_req
      -- CP-element group 356: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_word_addrgen/root_register_ack
      -- 
    ack_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1095_delayed_8_0_1101_inst_ack_1, ack => maxPool4_CP_360_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	87 
    -- CP-element group 357: 	91 
    -- CP-element group 357: 	95 
    -- CP-element group 357: 	99 
    -- CP-element group 357: 	151 
    -- CP-element group 357: 	155 
    -- CP-element group 357: 	159 
    -- CP-element group 357: 	163 
    -- CP-element group 357: 	215 
    -- CP-element group 357: 	219 
    -- CP-element group 357: 	223 
    -- CP-element group 357: 	227 
    -- CP-element group 357: 	279 
    -- CP-element group 357: 	283 
    -- CP-element group 357: 	287 
    -- CP-element group 357: 	291 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_sample_start_
      -- CP-element group 357: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Sample/$entry
      -- CP-element group 357: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Sample/rr
      -- 
    rr_1973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(357), ack => CONCAT_u32_u64_1116_inst_req_0); -- 
    maxPool4_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(87) & maxPool4_CP_360_elements(91) & maxPool4_CP_360_elements(95) & maxPool4_CP_360_elements(99) & maxPool4_CP_360_elements(151) & maxPool4_CP_360_elements(155) & maxPool4_CP_360_elements(159) & maxPool4_CP_360_elements(163) & maxPool4_CP_360_elements(215) & maxPool4_CP_360_elements(219) & maxPool4_CP_360_elements(223) & maxPool4_CP_360_elements(227) & maxPool4_CP_360_elements(279) & maxPool4_CP_360_elements(283) & maxPool4_CP_360_elements(287) & maxPool4_CP_360_elements(291) & maxPool4_CP_360_elements(359);
      gj_maxPool4_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: 	363 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_update_start_
      -- CP-element group 358: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Update/$entry
      -- CP-element group 358: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Update/cr
      -- 
    cr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(358), ack => CONCAT_u32_u64_1116_inst_req_1); -- 
    maxPool4_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(360) & maxPool4_CP_360_elements(363);
      gj_maxPool4_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	85 
    -- CP-element group 359: 	89 
    -- CP-element group 359: 	93 
    -- CP-element group 359: 	97 
    -- CP-element group 359: 	149 
    -- CP-element group 359: 	153 
    -- CP-element group 359: 	157 
    -- CP-element group 359: 	161 
    -- CP-element group 359: 	213 
    -- CP-element group 359: 	217 
    -- CP-element group 359: 	221 
    -- CP-element group 359: 	225 
    -- CP-element group 359: 	277 
    -- CP-element group 359: 	281 
    -- CP-element group 359: 	285 
    -- CP-element group 359: 	289 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_sample_completed_
      -- CP-element group 359: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Sample/$exit
      -- CP-element group 359: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Sample/ra
      -- 
    ra_1974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1116_inst_ack_0, ack => maxPool4_CP_360_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_update_completed_
      -- CP-element group 360: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Update/$exit
      -- CP-element group 360: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1116_Update/ca
      -- 
    ca_1979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1116_inst_ack_1, ack => maxPool4_CP_360_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	356 
    -- CP-element group 361: 	360 
    -- CP-element group 361: 	389 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (9) 
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_sample_start_
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/$entry
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/ptr_deref_1105_Split/$entry
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/ptr_deref_1105_Split/$exit
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/ptr_deref_1105_Split/split_req
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/ptr_deref_1105_Split/split_ack
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/$entry
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/word_0/$entry
      -- CP-element group 361: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/word_0/rr
      -- 
    rr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(361), ack => ptr_deref_1105_store_0_req_0); -- 
    maxPool4_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(356) & maxPool4_CP_360_elements(360) & maxPool4_CP_360_elements(389) & maxPool4_CP_360_elements(363);
      gj_maxPool4_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_update_start_
      -- CP-element group 362: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/$entry
      -- CP-element group 362: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/$entry
      -- CP-element group 362: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/word_0/$entry
      -- CP-element group 362: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/word_0/cr
      -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(362), ack => ptr_deref_1105_store_0_req_1); -- 
    maxPool4_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(364);
      gj_maxPool4_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	390 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	354 
    -- CP-element group 363: 	358 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_sample_completed_
      -- CP-element group 363: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/$exit
      -- CP-element group 363: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/$exit
      -- CP-element group 363: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/word_0/$exit
      -- CP-element group 363: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Sample/word_access_start/word_0/ra
      -- 
    ra_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_store_0_ack_0, ack => maxPool4_CP_360_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	391 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_update_completed_
      -- CP-element group 364: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/$exit
      -- CP-element group 364: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/$exit
      -- CP-element group 364: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/word_0/$exit
      -- CP-element group 364: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_Update/word_access_complete/word_0/ca
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1105_store_0_ack_1, ack => maxPool4_CP_360_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	369 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	370 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	370 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_sample_start_
      -- CP-element group 365: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_request/$entry
      -- CP-element group 365: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_request/req
      -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(365), ack => addr_of_1125_final_reg_req_0); -- 
    maxPool4_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(369) & maxPool4_CP_360_elements(370);
      gj_maxPool4_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	1 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	371 
    -- CP-element group 366: 	374 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	371 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_update_start_
      -- CP-element group 366: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_complete/$entry
      -- CP-element group 366: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_complete/req
      -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(366), ack => addr_of_1125_final_reg_req_1); -- 
    maxPool4_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(371) & maxPool4_CP_360_elements(374);
      gj_maxPool4_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	1 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: 	370 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_update_start
      -- CP-element group 367: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Update/$entry
      -- CP-element group 367: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Update/req
      -- 
    req_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(367), ack => array_obj_ref_1124_index_offset_req_1); -- 
    maxPool4_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(1) & maxPool4_CP_360_elements(369) & maxPool4_CP_360_elements(370);
      gj_maxPool4_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	1 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	391 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	2 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_sample_complete
      -- CP-element group 368: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Sample/$exit
      -- CP-element group 368: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Sample/ack
      -- 
    ack_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1124_index_offset_ack_0, ack => maxPool4_CP_360_elements(368)); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (8) 
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_root_address_calculated
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_offset_calculated
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Update/$exit
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_final_index_sum_regn_Update/ack
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_base_plus_offset/$entry
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_base_plus_offset/$exit
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 assign_stmt_106_to_assign_stmt_1147/array_obj_ref_1124_base_plus_offset/sum_rename_ack
      -- 
    ack_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1124_index_offset_ack_1, ack => maxPool4_CP_360_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: 	367 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_sample_completed_
      -- CP-element group 370: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_request/$exit
      -- CP-element group 370: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_request/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1125_final_reg_ack_0, ack => maxPool4_CP_360_elements(370)); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	366 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	366 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_update_completed_
      -- CP-element group 371: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_complete/$exit
      -- CP-element group 371: 	 assign_stmt_106_to_assign_stmt_1147/addr_of_1125_complete/ack
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1125_final_reg_ack_1, ack => maxPool4_CP_360_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_sample_start_
      -- CP-element group 372: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Sample/$entry
      -- CP-element group 372: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Sample/req
      -- 
    req_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(372), ack => W_myptr8_1118_delayed_8_0_1127_inst_req_0); -- 
    maxPool4_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(371) & maxPool4_CP_360_elements(374);
      gj_maxPool4_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	382 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_update_start_
      -- CP-element group 373: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Update/$entry
      -- CP-element group 373: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Update/req
      -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(373), ack => W_myptr8_1118_delayed_8_0_1127_inst_req_1); -- 
    maxPool4_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(375) & maxPool4_CP_360_elements(382);
      gj_maxPool4_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_sample_completed_
      -- CP-element group 374: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Sample/$exit
      -- CP-element group 374: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Sample/ack
      -- 
    ack_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1118_delayed_8_0_1127_inst_ack_0, ack => maxPool4_CP_360_elements(374)); -- 
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	380 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (19) 
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_update_completed_
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Update/$exit
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/assign_stmt_1129_Update/ack
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_address_calculated
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_word_address_calculated
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_root_address_calculated
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_address_resized
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_addr_resize/$entry
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_addr_resize/$exit
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_addr_resize/base_resize_req
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_addr_resize/base_resize_ack
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_plus_offset/$entry
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_plus_offset/$exit
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_plus_offset/sum_rename_req
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_base_plus_offset/sum_rename_ack
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_word_addrgen/$entry
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_word_addrgen/$exit
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_word_addrgen/root_register_req
      -- CP-element group 375: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_word_addrgen/root_register_ack
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1118_delayed_8_0_1127_inst_ack_1, ack => maxPool4_CP_360_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	103 
    -- CP-element group 376: 	107 
    -- CP-element group 376: 	111 
    -- CP-element group 376: 	115 
    -- CP-element group 376: 	167 
    -- CP-element group 376: 	171 
    -- CP-element group 376: 	175 
    -- CP-element group 376: 	179 
    -- CP-element group 376: 	231 
    -- CP-element group 376: 	235 
    -- CP-element group 376: 	239 
    -- CP-element group 376: 	243 
    -- CP-element group 376: 	295 
    -- CP-element group 376: 	299 
    -- CP-element group 376: 	303 
    -- CP-element group 376: 	307 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_sample_start_
      -- CP-element group 376: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Sample/$entry
      -- CP-element group 376: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Sample/rr
      -- 
    rr_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(376), ack => CONCAT_u32_u64_1142_inst_req_0); -- 
    maxPool4_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(103) & maxPool4_CP_360_elements(107) & maxPool4_CP_360_elements(111) & maxPool4_CP_360_elements(115) & maxPool4_CP_360_elements(167) & maxPool4_CP_360_elements(171) & maxPool4_CP_360_elements(175) & maxPool4_CP_360_elements(179) & maxPool4_CP_360_elements(231) & maxPool4_CP_360_elements(235) & maxPool4_CP_360_elements(239) & maxPool4_CP_360_elements(243) & maxPool4_CP_360_elements(295) & maxPool4_CP_360_elements(299) & maxPool4_CP_360_elements(303) & maxPool4_CP_360_elements(307) & maxPool4_CP_360_elements(378);
      gj_maxPool4_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: 	382 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_update_start_
      -- CP-element group 377: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Update/$entry
      -- CP-element group 377: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Update/cr
      -- 
    cr_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(377), ack => CONCAT_u32_u64_1142_inst_req_1); -- 
    maxPool4_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(379) & maxPool4_CP_360_elements(382);
      gj_maxPool4_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	101 
    -- CP-element group 378: 	105 
    -- CP-element group 378: 	109 
    -- CP-element group 378: 	113 
    -- CP-element group 378: 	165 
    -- CP-element group 378: 	169 
    -- CP-element group 378: 	173 
    -- CP-element group 378: 	177 
    -- CP-element group 378: 	229 
    -- CP-element group 378: 	233 
    -- CP-element group 378: 	237 
    -- CP-element group 378: 	241 
    -- CP-element group 378: 	293 
    -- CP-element group 378: 	297 
    -- CP-element group 378: 	301 
    -- CP-element group 378: 	305 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_sample_completed_
      -- CP-element group 378: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Sample/$exit
      -- CP-element group 378: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Sample/ra
      -- 
    ra_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1142_inst_ack_0, ack => maxPool4_CP_360_elements(378)); -- 
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_update_completed_
      -- CP-element group 379: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Update/$exit
      -- CP-element group 379: 	 assign_stmt_106_to_assign_stmt_1147/CONCAT_u32_u64_1142_Update/ca
      -- 
    ca_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1142_inst_ack_1, ack => maxPool4_CP_360_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	375 
    -- CP-element group 380: 	379 
    -- CP-element group 380: 	390 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (9) 
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_sample_start_
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/$entry
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/ptr_deref_1131_Split/$entry
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/ptr_deref_1131_Split/$exit
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/ptr_deref_1131_Split/split_req
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/ptr_deref_1131_Split/split_ack
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/$entry
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/word_0/rr
      -- 
    rr_2141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(380), ack => ptr_deref_1131_store_0_req_0); -- 
    maxPool4_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(375) & maxPool4_CP_360_elements(379) & maxPool4_CP_360_elements(390) & maxPool4_CP_360_elements(382);
      gj_maxPool4_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_update_start_
      -- CP-element group 381: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/$entry
      -- CP-element group 381: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/$entry
      -- CP-element group 381: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/word_0/$entry
      -- CP-element group 381: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/word_0/cr
      -- 
    cr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(381), ack => ptr_deref_1131_store_0_req_1); -- 
    maxPool4_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_360_elements(383);
      gj_maxPool4_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	391 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	323 
    -- CP-element group 382: 	373 
    -- CP-element group 382: 	377 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_sample_completed_
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/$exit
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/$exit
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/word_0/$exit
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Sample/word_access_start/word_0/ra
      -- CP-element group 382: 	 assign_stmt_106_to_assign_stmt_1147/ring_reenable_memory_space_0
      -- 
    ra_2142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1131_store_0_ack_0, ack => maxPool4_CP_360_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	391 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_update_completed_
      -- CP-element group 383: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/$exit
      -- CP-element group 383: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/$exit
      -- CP-element group 383: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/word_0/$exit
      -- CP-element group 383: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1131_Update/word_access_complete/word_0/ca
      -- 
    ca_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1131_store_0_ack_1, ack => maxPool4_CP_360_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	55 
    -- CP-element group 384: 	119 
    -- CP-element group 384: 	183 
    -- CP-element group 384: 	247 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_sample_start_
      -- CP-element group 384: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Sample/$entry
      -- CP-element group 384: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Sample/rr
      -- 
    rr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(384), ack => type_cast_1146_inst_req_0); -- 
    maxPool4_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(55) & maxPool4_CP_360_elements(119) & maxPool4_CP_360_elements(183) & maxPool4_CP_360_elements(247) & maxPool4_CP_360_elements(386);
      gj_maxPool4_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	7 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_update_start_
      -- CP-element group 385: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Update/$entry
      -- CP-element group 385: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Update/cr
      -- 
    cr_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_360_elements(385), ack => type_cast_1146_inst_req_1); -- 
    maxPool4_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(7) & maxPool4_CP_360_elements(387);
      gj_maxPool4_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	53 
    -- CP-element group 386: 	117 
    -- CP-element group 386: 	181 
    -- CP-element group 386: 	245 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_sample_completed_
      -- CP-element group 386: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Sample/$exit
      -- CP-element group 386: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Sample/ra
      -- 
    ra_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1146_inst_ack_0, ack => maxPool4_CP_360_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	391 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_update_completed_
      -- CP-element group 387: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Update/$exit
      -- CP-element group 387: 	 assign_stmt_106_to_assign_stmt_1147/type_cast_1146_Update/ca
      -- 
    ca_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1146_inst_ack_1, ack => maxPool4_CP_360_elements(387)); -- 
    -- CP-element group 388:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	325 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	342 
    -- CP-element group 388:  members (1) 
      -- CP-element group 388: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1053_ptr_deref_1079_delay
      -- 
    -- Element group maxPool4_CP_360_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => maxPool4_CP_360_elements(325), ack => maxPool4_CP_360_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	344 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	361 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1079_ptr_deref_1105_delay
      -- 
    -- Element group maxPool4_CP_360_elements(389) is a control-delay.
    cp_element_389_delay: control_delay_element  generic map(name => " 389_delay", delay_value => 1)  port map(req => maxPool4_CP_360_elements(344), ack => maxPool4_CP_360_elements(389), clk => clk, reset =>reset);
    -- CP-element group 390:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	363 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	380 
    -- CP-element group 390:  members (1) 
      -- CP-element group 390: 	 assign_stmt_106_to_assign_stmt_1147/ptr_deref_1105_ptr_deref_1131_delay
      -- 
    -- Element group maxPool4_CP_360_elements(390) is a control-delay.
    cp_element_390_delay: control_delay_element  generic map(name => " 390_delay", delay_value => 1)  port map(req => maxPool4_CP_360_elements(363), ack => maxPool4_CP_360_elements(390), clk => clk, reset =>reset);
    -- CP-element group 391:  join  transition  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	11 
    -- CP-element group 391: 	18 
    -- CP-element group 391: 	25 
    -- CP-element group 391: 	32 
    -- CP-element group 391: 	311 
    -- CP-element group 391: 	326 
    -- CP-element group 391: 	330 
    -- CP-element group 391: 	345 
    -- CP-element group 391: 	349 
    -- CP-element group 391: 	364 
    -- CP-element group 391: 	368 
    -- CP-element group 391: 	382 
    -- CP-element group 391: 	383 
    -- CP-element group 391: 	387 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	398 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 assign_stmt_106_to_assign_stmt_1147/$exit
      -- 
    maxPool4_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= maxPool4_CP_360_elements(11) & maxPool4_CP_360_elements(18) & maxPool4_CP_360_elements(25) & maxPool4_CP_360_elements(32) & maxPool4_CP_360_elements(311) & maxPool4_CP_360_elements(326) & maxPool4_CP_360_elements(330) & maxPool4_CP_360_elements(345) & maxPool4_CP_360_elements(349) & maxPool4_CP_360_elements(364) & maxPool4_CP_360_elements(368) & maxPool4_CP_360_elements(382) & maxPool4_CP_360_elements(383) & maxPool4_CP_360_elements(387);
      gj_maxPool4_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_360_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  place  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	2 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 addr_update_enable
      -- 
    maxPool4_CP_360_elements(392) <= maxPool4_CP_360_elements(2);
    -- CP-element group 393:  place  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	3 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 addr1_update_enable
      -- 
    maxPool4_CP_360_elements(393) <= maxPool4_CP_360_elements(3);
    -- CP-element group 394:  place  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	4 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 addr2_update_enable
      -- 
    maxPool4_CP_360_elements(394) <= maxPool4_CP_360_elements(4);
    -- CP-element group 395:  place  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	5 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 addr3_update_enable
      -- 
    maxPool4_CP_360_elements(395) <= maxPool4_CP_360_elements(5);
    -- CP-element group 396:  place  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	6 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 addr4_update_enable
      -- 
    maxPool4_CP_360_elements(396) <= maxPool4_CP_360_elements(6);
    -- CP-element group 397:  place  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	7 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 output_update_enable
      -- 
    -- CP-element group 398:  transition  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	391 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (1) 
      -- CP-element group 398: 	 $exit
      -- 
    maxPool4_CP_360_elements(398) <= maxPool4_CP_360_elements(391);
    --  hookup: inputs to control-path 
    maxPool4_CP_360_elements(397) <= output_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= maxPool4_CP_360_elements(392);
    addr1_update_enable <= maxPool4_CP_360_elements(393);
    addr2_update_enable <= maxPool4_CP_360_elements(394);
    addr3_update_enable <= maxPool4_CP_360_elements(395);
    addr4_update_enable <= maxPool4_CP_360_elements(396);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1071_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1071_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1071_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1097_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1097_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1097_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1123_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1123_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1123_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1058_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1063_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1084_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1089_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1110_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1115_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1136_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1141_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_1064_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1090_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1116_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1142_wire : std_logic_vector(63 downto 0);
    signal R_addr1_103_resized : std_logic_vector(13 downto 0);
    signal R_addr1_103_scaled : std_logic_vector(13 downto 0);
    signal R_addr2_110_resized : std_logic_vector(13 downto 0);
    signal R_addr2_110_scaled : std_logic_vector(13 downto 0);
    signal R_addr3_117_resized : std_logic_vector(13 downto 0);
    signal R_addr3_117_scaled : std_logic_vector(13 downto 0);
    signal R_addr4_124_resized : std_logic_vector(13 downto 0);
    signal R_addr4_124_scaled : std_logic_vector(13 downto 0);
    signal R_addr_1045_resized : std_logic_vector(13 downto 0);
    signal R_addr_1045_scaled : std_logic_vector(13 downto 0);
    signal SGT_i16_u1_1005_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1013_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1021_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1029_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1037_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_661_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_669_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_677_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_685_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_693_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_701_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_709_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_717_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_725_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_733_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_741_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_749_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_757_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_765_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_773_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_781_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_789_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_797_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_805_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_813_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_821_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_829_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_837_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_845_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_853_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_861_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_869_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_877_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_885_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_893_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_901_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_909_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_917_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_925_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_933_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_941_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_949_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_957_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_965_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_973_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_981_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_989_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_997_wire : std_logic_vector(0 downto 0);
    signal a110_441 : std_logic_vector(15 downto 0);
    signal a111_445 : std_logic_vector(15 downto 0);
    signal a112_449 : std_logic_vector(15 downto 0);
    signal a113_453 : std_logic_vector(15 downto 0);
    signal a114_457 : std_logic_vector(15 downto 0);
    signal a115_461 : std_logic_vector(15 downto 0);
    signal a116_465 : std_logic_vector(15 downto 0);
    signal a11_405 : std_logic_vector(15 downto 0);
    signal a12_409 : std_logic_vector(15 downto 0);
    signal a13_413 : std_logic_vector(15 downto 0);
    signal a14_417 : std_logic_vector(15 downto 0);
    signal a15_421 : std_logic_vector(15 downto 0);
    signal a16_425 : std_logic_vector(15 downto 0);
    signal a17_429 : std_logic_vector(15 downto 0);
    signal a18_433 : std_logic_vector(15 downto 0);
    signal a19_437 : std_logic_vector(15 downto 0);
    signal a210_505 : std_logic_vector(15 downto 0);
    signal a211_509 : std_logic_vector(15 downto 0);
    signal a212_513 : std_logic_vector(15 downto 0);
    signal a213_517 : std_logic_vector(15 downto 0);
    signal a214_521 : std_logic_vector(15 downto 0);
    signal a215_525 : std_logic_vector(15 downto 0);
    signal a216_529 : std_logic_vector(15 downto 0);
    signal a21_469 : std_logic_vector(15 downto 0);
    signal a22_473 : std_logic_vector(15 downto 0);
    signal a23_477 : std_logic_vector(15 downto 0);
    signal a24_481 : std_logic_vector(15 downto 0);
    signal a25_485 : std_logic_vector(15 downto 0);
    signal a26_489 : std_logic_vector(15 downto 0);
    signal a27_493 : std_logic_vector(15 downto 0);
    signal a28_497 : std_logic_vector(15 downto 0);
    signal a29_501 : std_logic_vector(15 downto 0);
    signal a310_569 : std_logic_vector(15 downto 0);
    signal a311_573 : std_logic_vector(15 downto 0);
    signal a312_577 : std_logic_vector(15 downto 0);
    signal a313_581 : std_logic_vector(15 downto 0);
    signal a314_585 : std_logic_vector(15 downto 0);
    signal a315_589 : std_logic_vector(15 downto 0);
    signal a316_593 : std_logic_vector(15 downto 0);
    signal a31_533 : std_logic_vector(15 downto 0);
    signal a32_537 : std_logic_vector(15 downto 0);
    signal a33_541 : std_logic_vector(15 downto 0);
    signal a34_545 : std_logic_vector(15 downto 0);
    signal a35_549 : std_logic_vector(15 downto 0);
    signal a36_553 : std_logic_vector(15 downto 0);
    signal a37_557 : std_logic_vector(15 downto 0);
    signal a38_561 : std_logic_vector(15 downto 0);
    signal a39_565 : std_logic_vector(15 downto 0);
    signal a410_633 : std_logic_vector(15 downto 0);
    signal a411_637 : std_logic_vector(15 downto 0);
    signal a412_641 : std_logic_vector(15 downto 0);
    signal a413_645 : std_logic_vector(15 downto 0);
    signal a414_649 : std_logic_vector(15 downto 0);
    signal a415_653 : std_logic_vector(15 downto 0);
    signal a416_657 : std_logic_vector(15 downto 0);
    signal a41_597 : std_logic_vector(15 downto 0);
    signal a42_601 : std_logic_vector(15 downto 0);
    signal a43_605 : std_logic_vector(15 downto 0);
    signal a44_609 : std_logic_vector(15 downto 0);
    signal a45_613 : std_logic_vector(15 downto 0);
    signal a46_617 : std_logic_vector(15 downto 0);
    signal a47_621 : std_logic_vector(15 downto 0);
    signal a48_625 : std_logic_vector(15 downto 0);
    signal a49_629 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1046_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1046_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1046_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1046_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1046_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1046_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_104_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1072_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1098_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_111_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1124_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_118_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_125_root_address : std_logic_vector(13 downto 0);
    signal c1_131 : std_logic_vector(255 downto 0);
    signal c2_135 : std_logic_vector(255 downto 0);
    signal c3_139 : std_logic_vector(255 downto 0);
    signal c4_143 : std_logic_vector(255 downto 0);
    signal konst_1070_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1096_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1122_wire_constant : std_logic_vector(31 downto 0);
    signal myptr1_106 : std_logic_vector(31 downto 0);
    signal myptr2_113 : std_logic_vector(31 downto 0);
    signal myptr3_120 : std_logic_vector(31 downto 0);
    signal myptr4_127 : std_logic_vector(31 downto 0);
    signal myptr5_1048 : std_logic_vector(31 downto 0);
    signal myptr5_1049_delayed_8_0_1051 : std_logic_vector(31 downto 0);
    signal myptr6_1072_delayed_8_0_1077 : std_logic_vector(31 downto 0);
    signal myptr6_1074 : std_logic_vector(31 downto 0);
    signal myptr7_1095_delayed_8_0_1103 : std_logic_vector(31 downto 0);
    signal myptr7_1100 : std_logic_vector(31 downto 0);
    signal myptr8_1118_delayed_8_0_1129 : std_logic_vector(31 downto 0);
    signal myptr8_1126 : std_logic_vector(31 downto 0);
    signal out10_897 : std_logic_vector(15 downto 0);
    signal out11_921 : std_logic_vector(15 downto 0);
    signal out12_945 : std_logic_vector(15 downto 0);
    signal out13_969 : std_logic_vector(15 downto 0);
    signal out14_993 : std_logic_vector(15 downto 0);
    signal out15_1017 : std_logic_vector(15 downto 0);
    signal out16_1041 : std_logic_vector(15 downto 0);
    signal out1_681 : std_logic_vector(15 downto 0);
    signal out2_705 : std_logic_vector(15 downto 0);
    signal out3_729 : std_logic_vector(15 downto 0);
    signal out4_753 : std_logic_vector(15 downto 0);
    signal out5_777 : std_logic_vector(15 downto 0);
    signal out6_801 : std_logic_vector(15 downto 0);
    signal out7_825 : std_logic_vector(15 downto 0);
    signal out8_849 : std_logic_vector(15 downto 0);
    signal out9_873 : std_logic_vector(15 downto 0);
    signal ptr_deref_1053_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1053_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1053_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1053_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1053_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1053_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1079_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1079_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1079_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1079_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1079_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1079_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1105_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1105_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1105_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1105_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1105_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1105_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1131_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1131_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1131_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1131_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1131_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1131_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_130_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_130_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_130_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_130_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_130_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_134_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_134_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_134_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_134_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_134_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_142_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_142_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_142_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_142_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_142_word_offset_0 : std_logic_vector(13 downto 0);
    signal sliced_v110_184 : std_logic_vector(15 downto 0);
    signal sliced_v111_188 : std_logic_vector(15 downto 0);
    signal sliced_v112_192 : std_logic_vector(15 downto 0);
    signal sliced_v113_196 : std_logic_vector(15 downto 0);
    signal sliced_v114_200 : std_logic_vector(15 downto 0);
    signal sliced_v115_204 : std_logic_vector(15 downto 0);
    signal sliced_v116_208 : std_logic_vector(15 downto 0);
    signal sliced_v11_148 : std_logic_vector(15 downto 0);
    signal sliced_v12_152 : std_logic_vector(15 downto 0);
    signal sliced_v13_156 : std_logic_vector(15 downto 0);
    signal sliced_v14_160 : std_logic_vector(15 downto 0);
    signal sliced_v15_164 : std_logic_vector(15 downto 0);
    signal sliced_v16_168 : std_logic_vector(15 downto 0);
    signal sliced_v17_172 : std_logic_vector(15 downto 0);
    signal sliced_v18_176 : std_logic_vector(15 downto 0);
    signal sliced_v19_180 : std_logic_vector(15 downto 0);
    signal sliced_v210_248 : std_logic_vector(15 downto 0);
    signal sliced_v211_252 : std_logic_vector(15 downto 0);
    signal sliced_v212_256 : std_logic_vector(15 downto 0);
    signal sliced_v213_260 : std_logic_vector(15 downto 0);
    signal sliced_v214_264 : std_logic_vector(15 downto 0);
    signal sliced_v215_268 : std_logic_vector(15 downto 0);
    signal sliced_v216_272 : std_logic_vector(15 downto 0);
    signal sliced_v21_212 : std_logic_vector(15 downto 0);
    signal sliced_v22_216 : std_logic_vector(15 downto 0);
    signal sliced_v23_220 : std_logic_vector(15 downto 0);
    signal sliced_v24_224 : std_logic_vector(15 downto 0);
    signal sliced_v25_228 : std_logic_vector(15 downto 0);
    signal sliced_v26_232 : std_logic_vector(15 downto 0);
    signal sliced_v27_236 : std_logic_vector(15 downto 0);
    signal sliced_v28_240 : std_logic_vector(15 downto 0);
    signal sliced_v29_244 : std_logic_vector(15 downto 0);
    signal sliced_v310_312 : std_logic_vector(15 downto 0);
    signal sliced_v311_316 : std_logic_vector(15 downto 0);
    signal sliced_v312_320 : std_logic_vector(15 downto 0);
    signal sliced_v313_324 : std_logic_vector(15 downto 0);
    signal sliced_v314_328 : std_logic_vector(15 downto 0);
    signal sliced_v315_332 : std_logic_vector(15 downto 0);
    signal sliced_v316_336 : std_logic_vector(15 downto 0);
    signal sliced_v31_276 : std_logic_vector(15 downto 0);
    signal sliced_v32_280 : std_logic_vector(15 downto 0);
    signal sliced_v33_284 : std_logic_vector(15 downto 0);
    signal sliced_v34_288 : std_logic_vector(15 downto 0);
    signal sliced_v35_292 : std_logic_vector(15 downto 0);
    signal sliced_v36_296 : std_logic_vector(15 downto 0);
    signal sliced_v37_300 : std_logic_vector(15 downto 0);
    signal sliced_v38_304 : std_logic_vector(15 downto 0);
    signal sliced_v39_308 : std_logic_vector(15 downto 0);
    signal sliced_v410_376 : std_logic_vector(15 downto 0);
    signal sliced_v411_380 : std_logic_vector(15 downto 0);
    signal sliced_v412_384 : std_logic_vector(15 downto 0);
    signal sliced_v413_388 : std_logic_vector(15 downto 0);
    signal sliced_v414_392 : std_logic_vector(15 downto 0);
    signal sliced_v415_396 : std_logic_vector(15 downto 0);
    signal sliced_v416_400 : std_logic_vector(15 downto 0);
    signal sliced_v41_340 : std_logic_vector(15 downto 0);
    signal sliced_v42_344 : std_logic_vector(15 downto 0);
    signal sliced_v43_348 : std_logic_vector(15 downto 0);
    signal sliced_v44_352 : std_logic_vector(15 downto 0);
    signal sliced_v45_356 : std_logic_vector(15 downto 0);
    signal sliced_v46_360 : std_logic_vector(15 downto 0);
    signal sliced_v47_364 : std_logic_vector(15 downto 0);
    signal sliced_v48_368 : std_logic_vector(15 downto 0);
    signal sliced_v49_372 : std_logic_vector(15 downto 0);
    signal t101_881 : std_logic_vector(15 downto 0);
    signal t102_889 : std_logic_vector(15 downto 0);
    signal t111_905 : std_logic_vector(15 downto 0);
    signal t112_913 : std_logic_vector(15 downto 0);
    signal t11_665 : std_logic_vector(15 downto 0);
    signal t121_929 : std_logic_vector(15 downto 0);
    signal t122_937 : std_logic_vector(15 downto 0);
    signal t12_673 : std_logic_vector(15 downto 0);
    signal t131_953 : std_logic_vector(15 downto 0);
    signal t132_961 : std_logic_vector(15 downto 0);
    signal t141_977 : std_logic_vector(15 downto 0);
    signal t142_985 : std_logic_vector(15 downto 0);
    signal t151_1001 : std_logic_vector(15 downto 0);
    signal t152_1009 : std_logic_vector(15 downto 0);
    signal t161_1025 : std_logic_vector(15 downto 0);
    signal t162_1033 : std_logic_vector(15 downto 0);
    signal t21_689 : std_logic_vector(15 downto 0);
    signal t22_697 : std_logic_vector(15 downto 0);
    signal t31_713 : std_logic_vector(15 downto 0);
    signal t32_721 : std_logic_vector(15 downto 0);
    signal t41_737 : std_logic_vector(15 downto 0);
    signal t42_745 : std_logic_vector(15 downto 0);
    signal t51_761 : std_logic_vector(15 downto 0);
    signal t52_769 : std_logic_vector(15 downto 0);
    signal t61_785 : std_logic_vector(15 downto 0);
    signal t62_793 : std_logic_vector(15 downto 0);
    signal t71_809 : std_logic_vector(15 downto 0);
    signal t72_817 : std_logic_vector(15 downto 0);
    signal t81_833 : std_logic_vector(15 downto 0);
    signal t82_841 : std_logic_vector(15 downto 0);
    signal t91_857 : std_logic_vector(15 downto 0);
    signal t92_865 : std_logic_vector(15 downto 0);
    signal type_cast_1055_wire : std_logic_vector(15 downto 0);
    signal type_cast_1057_wire : std_logic_vector(15 downto 0);
    signal type_cast_1060_wire : std_logic_vector(15 downto 0);
    signal type_cast_1062_wire : std_logic_vector(15 downto 0);
    signal type_cast_1081_wire : std_logic_vector(15 downto 0);
    signal type_cast_1083_wire : std_logic_vector(15 downto 0);
    signal type_cast_1086_wire : std_logic_vector(15 downto 0);
    signal type_cast_1088_wire : std_logic_vector(15 downto 0);
    signal type_cast_1107_wire : std_logic_vector(15 downto 0);
    signal type_cast_1109_wire : std_logic_vector(15 downto 0);
    signal type_cast_1112_wire : std_logic_vector(15 downto 0);
    signal type_cast_1114_wire : std_logic_vector(15 downto 0);
    signal type_cast_1133_wire : std_logic_vector(15 downto 0);
    signal type_cast_1135_wire : std_logic_vector(15 downto 0);
    signal type_cast_1138_wire : std_logic_vector(15 downto 0);
    signal type_cast_1140_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1046_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1046_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1046_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1046_resized_base_address <= "00000000000000";
    array_obj_ref_104_constant_part_of_offset <= "00000000000000";
    array_obj_ref_104_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_104_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_104_resized_base_address <= "00000000000000";
    array_obj_ref_1072_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1072_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1072_resized_base_address <= "00000000000000";
    array_obj_ref_1098_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1098_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1098_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1098_resized_base_address <= "00000000000000";
    array_obj_ref_111_constant_part_of_offset <= "00000000000000";
    array_obj_ref_111_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_111_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_111_resized_base_address <= "00000000000000";
    array_obj_ref_1124_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1124_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1124_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1124_resized_base_address <= "00000000000000";
    array_obj_ref_118_constant_part_of_offset <= "00000000000000";
    array_obj_ref_118_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_118_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_118_resized_base_address <= "00000000000000";
    array_obj_ref_125_constant_part_of_offset <= "00000000000000";
    array_obj_ref_125_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_125_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_125_resized_base_address <= "00000000000000";
    konst_1070_wire_constant <= "00000000000000000000000000000001";
    konst_1096_wire_constant <= "00000000000000000000000000000010";
    konst_1122_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_1053_word_offset_0 <= "00000000000000";
    ptr_deref_1079_word_offset_0 <= "00000000000000";
    ptr_deref_1105_word_offset_0 <= "00000000000000";
    ptr_deref_1131_word_offset_0 <= "00000000000000";
    ptr_deref_130_word_offset_0 <= "00000000000000";
    ptr_deref_134_word_offset_0 <= "00000000000000";
    ptr_deref_138_word_offset_0 <= "00000000000000";
    ptr_deref_142_word_offset_0 <= "00000000000000";
    -- flow-through select operator MUX_1000_inst
    t151_1001 <= a115_461 when (SGT_i16_u1_997_wire(0) /=  '0') else a215_525;
    -- flow-through select operator MUX_1008_inst
    t152_1009 <= a315_589 when (SGT_i16_u1_1005_wire(0) /=  '0') else a415_653;
    -- flow-through select operator MUX_1016_inst
    out15_1017 <= t151_1001 when (SGT_i16_u1_1013_wire(0) /=  '0') else t152_1009;
    -- flow-through select operator MUX_1024_inst
    t161_1025 <= a116_465 when (SGT_i16_u1_1021_wire(0) /=  '0') else a216_529;
    -- flow-through select operator MUX_1032_inst
    t162_1033 <= a316_593 when (SGT_i16_u1_1029_wire(0) /=  '0') else a416_657;
    -- flow-through select operator MUX_1040_inst
    out16_1041 <= t161_1025 when (SGT_i16_u1_1037_wire(0) /=  '0') else t162_1033;
    -- flow-through select operator MUX_664_inst
    t11_665 <= a11_405 when (SGT_i16_u1_661_wire(0) /=  '0') else a21_469;
    -- flow-through select operator MUX_672_inst
    t12_673 <= a31_533 when (SGT_i16_u1_669_wire(0) /=  '0') else a41_597;
    -- flow-through select operator MUX_680_inst
    out1_681 <= t11_665 when (SGT_i16_u1_677_wire(0) /=  '0') else t12_673;
    -- flow-through select operator MUX_688_inst
    t21_689 <= a12_409 when (SGT_i16_u1_685_wire(0) /=  '0') else a22_473;
    -- flow-through select operator MUX_696_inst
    t22_697 <= a32_537 when (SGT_i16_u1_693_wire(0) /=  '0') else a42_601;
    -- flow-through select operator MUX_704_inst
    out2_705 <= t21_689 when (SGT_i16_u1_701_wire(0) /=  '0') else t22_697;
    -- flow-through select operator MUX_712_inst
    t31_713 <= a13_413 when (SGT_i16_u1_709_wire(0) /=  '0') else a23_477;
    -- flow-through select operator MUX_720_inst
    t32_721 <= a33_541 when (SGT_i16_u1_717_wire(0) /=  '0') else a43_605;
    -- flow-through select operator MUX_728_inst
    out3_729 <= t31_713 when (SGT_i16_u1_725_wire(0) /=  '0') else t32_721;
    -- flow-through select operator MUX_736_inst
    t41_737 <= a14_417 when (SGT_i16_u1_733_wire(0) /=  '0') else a24_481;
    -- flow-through select operator MUX_744_inst
    t42_745 <= a34_545 when (SGT_i16_u1_741_wire(0) /=  '0') else a44_609;
    -- flow-through select operator MUX_752_inst
    out4_753 <= t41_737 when (SGT_i16_u1_749_wire(0) /=  '0') else t42_745;
    -- flow-through select operator MUX_760_inst
    t51_761 <= a15_421 when (SGT_i16_u1_757_wire(0) /=  '0') else a25_485;
    -- flow-through select operator MUX_768_inst
    t52_769 <= a35_549 when (SGT_i16_u1_765_wire(0) /=  '0') else a45_613;
    -- flow-through select operator MUX_776_inst
    out5_777 <= t51_761 when (SGT_i16_u1_773_wire(0) /=  '0') else t52_769;
    -- flow-through select operator MUX_784_inst
    t61_785 <= a16_425 when (SGT_i16_u1_781_wire(0) /=  '0') else a26_489;
    -- flow-through select operator MUX_792_inst
    t62_793 <= a36_553 when (SGT_i16_u1_789_wire(0) /=  '0') else a46_617;
    -- flow-through select operator MUX_800_inst
    out6_801 <= t61_785 when (SGT_i16_u1_797_wire(0) /=  '0') else t62_793;
    -- flow-through select operator MUX_808_inst
    t71_809 <= a17_429 when (SGT_i16_u1_805_wire(0) /=  '0') else a27_493;
    -- flow-through select operator MUX_816_inst
    t72_817 <= a37_557 when (SGT_i16_u1_813_wire(0) /=  '0') else a47_621;
    -- flow-through select operator MUX_824_inst
    out7_825 <= t71_809 when (SGT_i16_u1_821_wire(0) /=  '0') else t72_817;
    -- flow-through select operator MUX_832_inst
    t81_833 <= a18_433 when (SGT_i16_u1_829_wire(0) /=  '0') else a28_497;
    -- flow-through select operator MUX_840_inst
    t82_841 <= a38_561 when (SGT_i16_u1_837_wire(0) /=  '0') else a48_625;
    -- flow-through select operator MUX_848_inst
    out8_849 <= t81_833 when (SGT_i16_u1_845_wire(0) /=  '0') else t82_841;
    -- flow-through select operator MUX_856_inst
    t91_857 <= a19_437 when (SGT_i16_u1_853_wire(0) /=  '0') else a29_501;
    -- flow-through select operator MUX_864_inst
    t92_865 <= a39_565 when (SGT_i16_u1_861_wire(0) /=  '0') else a49_629;
    -- flow-through select operator MUX_872_inst
    out9_873 <= t91_857 when (SGT_i16_u1_869_wire(0) /=  '0') else t92_865;
    -- flow-through select operator MUX_880_inst
    t101_881 <= a110_441 when (SGT_i16_u1_877_wire(0) /=  '0') else a210_505;
    -- flow-through select operator MUX_888_inst
    t102_889 <= a310_569 when (SGT_i16_u1_885_wire(0) /=  '0') else a410_633;
    -- flow-through select operator MUX_896_inst
    out10_897 <= t101_881 when (SGT_i16_u1_893_wire(0) /=  '0') else t102_889;
    -- flow-through select operator MUX_904_inst
    t111_905 <= a111_445 when (SGT_i16_u1_901_wire(0) /=  '0') else a211_509;
    -- flow-through select operator MUX_912_inst
    t112_913 <= a311_573 when (SGT_i16_u1_909_wire(0) /=  '0') else a411_637;
    -- flow-through select operator MUX_920_inst
    out11_921 <= t111_905 when (SGT_i16_u1_917_wire(0) /=  '0') else t112_913;
    -- flow-through select operator MUX_928_inst
    t121_929 <= a112_449 when (SGT_i16_u1_925_wire(0) /=  '0') else a212_513;
    -- flow-through select operator MUX_936_inst
    t122_937 <= a312_577 when (SGT_i16_u1_933_wire(0) /=  '0') else a412_641;
    -- flow-through select operator MUX_944_inst
    out12_945 <= t121_929 when (SGT_i16_u1_941_wire(0) /=  '0') else t122_937;
    -- flow-through select operator MUX_952_inst
    t131_953 <= a113_453 when (SGT_i16_u1_949_wire(0) /=  '0') else a213_517;
    -- flow-through select operator MUX_960_inst
    t132_961 <= a313_581 when (SGT_i16_u1_957_wire(0) /=  '0') else a413_645;
    -- flow-through select operator MUX_968_inst
    out13_969 <= t131_953 when (SGT_i16_u1_965_wire(0) /=  '0') else t132_961;
    -- flow-through select operator MUX_976_inst
    t141_977 <= a114_457 when (SGT_i16_u1_973_wire(0) /=  '0') else a214_521;
    -- flow-through select operator MUX_984_inst
    t142_985 <= a314_585 when (SGT_i16_u1_981_wire(0) /=  '0') else a414_649;
    -- flow-through select operator MUX_992_inst
    out14_993 <= t141_977 when (SGT_i16_u1_989_wire(0) /=  '0') else t142_985;
    slice_147_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_147_inst_req_0;
      slice_147_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_147_inst_req_1;
      slice_147_inst_ack_1<= update_ack(0);
      slice_147_inst: SliceSplitProtocol generic map(name => "slice_147_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v11_148, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_151_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_151_inst_req_0;
      slice_151_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_151_inst_req_1;
      slice_151_inst_ack_1<= update_ack(0);
      slice_151_inst: SliceSplitProtocol generic map(name => "slice_151_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v12_152, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_155_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_155_inst_req_0;
      slice_155_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_155_inst_req_1;
      slice_155_inst_ack_1<= update_ack(0);
      slice_155_inst: SliceSplitProtocol generic map(name => "slice_155_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v13_156, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_159_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_159_inst_req_0;
      slice_159_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_159_inst_req_1;
      slice_159_inst_ack_1<= update_ack(0);
      slice_159_inst: SliceSplitProtocol generic map(name => "slice_159_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v14_160, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_163_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_163_inst_req_0;
      slice_163_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_163_inst_req_1;
      slice_163_inst_ack_1<= update_ack(0);
      slice_163_inst: SliceSplitProtocol generic map(name => "slice_163_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v15_164, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_167_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_167_inst_req_0;
      slice_167_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_167_inst_req_1;
      slice_167_inst_ack_1<= update_ack(0);
      slice_167_inst: SliceSplitProtocol generic map(name => "slice_167_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v16_168, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_171_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_171_inst_req_0;
      slice_171_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_171_inst_req_1;
      slice_171_inst_ack_1<= update_ack(0);
      slice_171_inst: SliceSplitProtocol generic map(name => "slice_171_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v17_172, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_175_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_175_inst_req_0;
      slice_175_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_175_inst_req_1;
      slice_175_inst_ack_1<= update_ack(0);
      slice_175_inst: SliceSplitProtocol generic map(name => "slice_175_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v18_176, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_179_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_179_inst_req_0;
      slice_179_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_179_inst_req_1;
      slice_179_inst_ack_1<= update_ack(0);
      slice_179_inst: SliceSplitProtocol generic map(name => "slice_179_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v19_180, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_183_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_183_inst_req_0;
      slice_183_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_183_inst_req_1;
      slice_183_inst_ack_1<= update_ack(0);
      slice_183_inst: SliceSplitProtocol generic map(name => "slice_183_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v110_184, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_187_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_187_inst_req_0;
      slice_187_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_187_inst_req_1;
      slice_187_inst_ack_1<= update_ack(0);
      slice_187_inst: SliceSplitProtocol generic map(name => "slice_187_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v111_188, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_191_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_191_inst_req_0;
      slice_191_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_191_inst_req_1;
      slice_191_inst_ack_1<= update_ack(0);
      slice_191_inst: SliceSplitProtocol generic map(name => "slice_191_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v112_192, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_195_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_195_inst_req_0;
      slice_195_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_195_inst_req_1;
      slice_195_inst_ack_1<= update_ack(0);
      slice_195_inst: SliceSplitProtocol generic map(name => "slice_195_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v113_196, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_199_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_199_inst_req_0;
      slice_199_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_199_inst_req_1;
      slice_199_inst_ack_1<= update_ack(0);
      slice_199_inst: SliceSplitProtocol generic map(name => "slice_199_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v114_200, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_203_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_203_inst_req_0;
      slice_203_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_203_inst_req_1;
      slice_203_inst_ack_1<= update_ack(0);
      slice_203_inst: SliceSplitProtocol generic map(name => "slice_203_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v115_204, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_207_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_207_inst_req_0;
      slice_207_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_207_inst_req_1;
      slice_207_inst_ack_1<= update_ack(0);
      slice_207_inst: SliceSplitProtocol generic map(name => "slice_207_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_131, dout => sliced_v116_208, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_211_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_211_inst_req_0;
      slice_211_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_211_inst_req_1;
      slice_211_inst_ack_1<= update_ack(0);
      slice_211_inst: SliceSplitProtocol generic map(name => "slice_211_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v21_212, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_215_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_215_inst_req_0;
      slice_215_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_215_inst_req_1;
      slice_215_inst_ack_1<= update_ack(0);
      slice_215_inst: SliceSplitProtocol generic map(name => "slice_215_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v22_216, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_219_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_219_inst_req_0;
      slice_219_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_219_inst_req_1;
      slice_219_inst_ack_1<= update_ack(0);
      slice_219_inst: SliceSplitProtocol generic map(name => "slice_219_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v23_220, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_223_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_223_inst_req_0;
      slice_223_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_223_inst_req_1;
      slice_223_inst_ack_1<= update_ack(0);
      slice_223_inst: SliceSplitProtocol generic map(name => "slice_223_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v24_224, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_227_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_227_inst_req_0;
      slice_227_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_227_inst_req_1;
      slice_227_inst_ack_1<= update_ack(0);
      slice_227_inst: SliceSplitProtocol generic map(name => "slice_227_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v25_228, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_231_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_231_inst_req_0;
      slice_231_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_231_inst_req_1;
      slice_231_inst_ack_1<= update_ack(0);
      slice_231_inst: SliceSplitProtocol generic map(name => "slice_231_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v26_232, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_235_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_235_inst_req_0;
      slice_235_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_235_inst_req_1;
      slice_235_inst_ack_1<= update_ack(0);
      slice_235_inst: SliceSplitProtocol generic map(name => "slice_235_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v27_236, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_239_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_239_inst_req_0;
      slice_239_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_239_inst_req_1;
      slice_239_inst_ack_1<= update_ack(0);
      slice_239_inst: SliceSplitProtocol generic map(name => "slice_239_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v28_240, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_243_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_243_inst_req_0;
      slice_243_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_243_inst_req_1;
      slice_243_inst_ack_1<= update_ack(0);
      slice_243_inst: SliceSplitProtocol generic map(name => "slice_243_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v29_244, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_247_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_247_inst_req_0;
      slice_247_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_247_inst_req_1;
      slice_247_inst_ack_1<= update_ack(0);
      slice_247_inst: SliceSplitProtocol generic map(name => "slice_247_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v210_248, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_251_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_251_inst_req_0;
      slice_251_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_251_inst_req_1;
      slice_251_inst_ack_1<= update_ack(0);
      slice_251_inst: SliceSplitProtocol generic map(name => "slice_251_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v211_252, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_255_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_255_inst_req_0;
      slice_255_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_255_inst_req_1;
      slice_255_inst_ack_1<= update_ack(0);
      slice_255_inst: SliceSplitProtocol generic map(name => "slice_255_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v212_256, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_259_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_259_inst_req_0;
      slice_259_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_259_inst_req_1;
      slice_259_inst_ack_1<= update_ack(0);
      slice_259_inst: SliceSplitProtocol generic map(name => "slice_259_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v213_260, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_263_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_263_inst_req_0;
      slice_263_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_263_inst_req_1;
      slice_263_inst_ack_1<= update_ack(0);
      slice_263_inst: SliceSplitProtocol generic map(name => "slice_263_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v214_264, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_267_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_267_inst_req_0;
      slice_267_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_267_inst_req_1;
      slice_267_inst_ack_1<= update_ack(0);
      slice_267_inst: SliceSplitProtocol generic map(name => "slice_267_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v215_268, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_271_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_271_inst_req_0;
      slice_271_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_271_inst_req_1;
      slice_271_inst_ack_1<= update_ack(0);
      slice_271_inst: SliceSplitProtocol generic map(name => "slice_271_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_135, dout => sliced_v216_272, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_275_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_275_inst_req_0;
      slice_275_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_275_inst_req_1;
      slice_275_inst_ack_1<= update_ack(0);
      slice_275_inst: SliceSplitProtocol generic map(name => "slice_275_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v31_276, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_279_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_279_inst_req_0;
      slice_279_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_279_inst_req_1;
      slice_279_inst_ack_1<= update_ack(0);
      slice_279_inst: SliceSplitProtocol generic map(name => "slice_279_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v32_280, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_283_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_283_inst_req_0;
      slice_283_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_283_inst_req_1;
      slice_283_inst_ack_1<= update_ack(0);
      slice_283_inst: SliceSplitProtocol generic map(name => "slice_283_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v33_284, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_287_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_287_inst_req_0;
      slice_287_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_287_inst_req_1;
      slice_287_inst_ack_1<= update_ack(0);
      slice_287_inst: SliceSplitProtocol generic map(name => "slice_287_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v34_288, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_291_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_291_inst_req_0;
      slice_291_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_291_inst_req_1;
      slice_291_inst_ack_1<= update_ack(0);
      slice_291_inst: SliceSplitProtocol generic map(name => "slice_291_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v35_292, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_295_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_295_inst_req_0;
      slice_295_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_295_inst_req_1;
      slice_295_inst_ack_1<= update_ack(0);
      slice_295_inst: SliceSplitProtocol generic map(name => "slice_295_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v36_296, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_299_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_299_inst_req_0;
      slice_299_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_299_inst_req_1;
      slice_299_inst_ack_1<= update_ack(0);
      slice_299_inst: SliceSplitProtocol generic map(name => "slice_299_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v37_300, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_303_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_303_inst_req_0;
      slice_303_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_303_inst_req_1;
      slice_303_inst_ack_1<= update_ack(0);
      slice_303_inst: SliceSplitProtocol generic map(name => "slice_303_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v38_304, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_307_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_307_inst_req_0;
      slice_307_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_307_inst_req_1;
      slice_307_inst_ack_1<= update_ack(0);
      slice_307_inst: SliceSplitProtocol generic map(name => "slice_307_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v39_308, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_311_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_311_inst_req_0;
      slice_311_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_311_inst_req_1;
      slice_311_inst_ack_1<= update_ack(0);
      slice_311_inst: SliceSplitProtocol generic map(name => "slice_311_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v310_312, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_315_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_315_inst_req_0;
      slice_315_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_315_inst_req_1;
      slice_315_inst_ack_1<= update_ack(0);
      slice_315_inst: SliceSplitProtocol generic map(name => "slice_315_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v311_316, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_319_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_319_inst_req_0;
      slice_319_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_319_inst_req_1;
      slice_319_inst_ack_1<= update_ack(0);
      slice_319_inst: SliceSplitProtocol generic map(name => "slice_319_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v312_320, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_323_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_323_inst_req_0;
      slice_323_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_323_inst_req_1;
      slice_323_inst_ack_1<= update_ack(0);
      slice_323_inst: SliceSplitProtocol generic map(name => "slice_323_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v313_324, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_327_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_327_inst_req_0;
      slice_327_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_327_inst_req_1;
      slice_327_inst_ack_1<= update_ack(0);
      slice_327_inst: SliceSplitProtocol generic map(name => "slice_327_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v314_328, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_331_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_331_inst_req_0;
      slice_331_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_331_inst_req_1;
      slice_331_inst_ack_1<= update_ack(0);
      slice_331_inst: SliceSplitProtocol generic map(name => "slice_331_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v315_332, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_335_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_335_inst_req_0;
      slice_335_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_335_inst_req_1;
      slice_335_inst_ack_1<= update_ack(0);
      slice_335_inst: SliceSplitProtocol generic map(name => "slice_335_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_139, dout => sliced_v316_336, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_339_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_339_inst_req_0;
      slice_339_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_339_inst_req_1;
      slice_339_inst_ack_1<= update_ack(0);
      slice_339_inst: SliceSplitProtocol generic map(name => "slice_339_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v41_340, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_343_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_343_inst_req_0;
      slice_343_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_343_inst_req_1;
      slice_343_inst_ack_1<= update_ack(0);
      slice_343_inst: SliceSplitProtocol generic map(name => "slice_343_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v42_344, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_347_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_347_inst_req_0;
      slice_347_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_347_inst_req_1;
      slice_347_inst_ack_1<= update_ack(0);
      slice_347_inst: SliceSplitProtocol generic map(name => "slice_347_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v43_348, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_351_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_351_inst_req_0;
      slice_351_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_351_inst_req_1;
      slice_351_inst_ack_1<= update_ack(0);
      slice_351_inst: SliceSplitProtocol generic map(name => "slice_351_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v44_352, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_355_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_355_inst_req_0;
      slice_355_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_355_inst_req_1;
      slice_355_inst_ack_1<= update_ack(0);
      slice_355_inst: SliceSplitProtocol generic map(name => "slice_355_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v45_356, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_359_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_359_inst_req_0;
      slice_359_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_359_inst_req_1;
      slice_359_inst_ack_1<= update_ack(0);
      slice_359_inst: SliceSplitProtocol generic map(name => "slice_359_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v46_360, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_363_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_363_inst_req_0;
      slice_363_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_363_inst_req_1;
      slice_363_inst_ack_1<= update_ack(0);
      slice_363_inst: SliceSplitProtocol generic map(name => "slice_363_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v47_364, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_367_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_367_inst_req_0;
      slice_367_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_367_inst_req_1;
      slice_367_inst_ack_1<= update_ack(0);
      slice_367_inst: SliceSplitProtocol generic map(name => "slice_367_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v48_368, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_371_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_371_inst_req_0;
      slice_371_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_371_inst_req_1;
      slice_371_inst_ack_1<= update_ack(0);
      slice_371_inst: SliceSplitProtocol generic map(name => "slice_371_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v49_372, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_375_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_375_inst_req_0;
      slice_375_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_375_inst_req_1;
      slice_375_inst_ack_1<= update_ack(0);
      slice_375_inst: SliceSplitProtocol generic map(name => "slice_375_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v410_376, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_379_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_379_inst_req_0;
      slice_379_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_379_inst_req_1;
      slice_379_inst_ack_1<= update_ack(0);
      slice_379_inst: SliceSplitProtocol generic map(name => "slice_379_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v411_380, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_383_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_383_inst_req_0;
      slice_383_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_383_inst_req_1;
      slice_383_inst_ack_1<= update_ack(0);
      slice_383_inst: SliceSplitProtocol generic map(name => "slice_383_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v412_384, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_387_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_387_inst_req_0;
      slice_387_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_387_inst_req_1;
      slice_387_inst_ack_1<= update_ack(0);
      slice_387_inst: SliceSplitProtocol generic map(name => "slice_387_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v413_388, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_391_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_391_inst_req_0;
      slice_391_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_391_inst_req_1;
      slice_391_inst_ack_1<= update_ack(0);
      slice_391_inst: SliceSplitProtocol generic map(name => "slice_391_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v414_392, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_395_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_395_inst_req_0;
      slice_395_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_395_inst_req_1;
      slice_395_inst_ack_1<= update_ack(0);
      slice_395_inst: SliceSplitProtocol generic map(name => "slice_395_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v415_396, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_399_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_399_inst_req_0;
      slice_399_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_399_inst_req_1;
      slice_399_inst_ack_1<= update_ack(0);
      slice_399_inst: SliceSplitProtocol generic map(name => "slice_399_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_143, dout => sliced_v416_400, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_myptr5_1049_delayed_8_0_1049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr5_1049_delayed_8_0_1049_inst_req_0;
      W_myptr5_1049_delayed_8_0_1049_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr5_1049_delayed_8_0_1049_inst_req_1;
      W_myptr5_1049_delayed_8_0_1049_inst_ack_1<= rack(0);
      W_myptr5_1049_delayed_8_0_1049_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr5_1049_delayed_8_0_1049_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr5_1048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1049_delayed_8_0_1051,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr6_1072_delayed_8_0_1075_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr6_1072_delayed_8_0_1075_inst_req_0;
      W_myptr6_1072_delayed_8_0_1075_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr6_1072_delayed_8_0_1075_inst_req_1;
      W_myptr6_1072_delayed_8_0_1075_inst_ack_1<= rack(0);
      W_myptr6_1072_delayed_8_0_1075_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr6_1072_delayed_8_0_1075_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr6_1074,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1072_delayed_8_0_1077,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr7_1095_delayed_8_0_1101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr7_1095_delayed_8_0_1101_inst_req_0;
      W_myptr7_1095_delayed_8_0_1101_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr7_1095_delayed_8_0_1101_inst_req_1;
      W_myptr7_1095_delayed_8_0_1101_inst_ack_1<= rack(0);
      W_myptr7_1095_delayed_8_0_1101_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr7_1095_delayed_8_0_1101_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr7_1100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1095_delayed_8_0_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr8_1118_delayed_8_0_1127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr8_1118_delayed_8_0_1127_inst_req_0;
      W_myptr8_1118_delayed_8_0_1127_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr8_1118_delayed_8_0_1127_inst_req_1;
      W_myptr8_1118_delayed_8_0_1127_inst_ack_1<= rack(0);
      W_myptr8_1118_delayed_8_0_1127_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr8_1118_delayed_8_0_1127_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr8_1126,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1118_delayed_8_0_1129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1047_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1047_final_reg_req_0;
      addr_of_1047_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1047_final_reg_req_1;
      addr_of_1047_final_reg_ack_1<= rack(0);
      addr_of_1047_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1047_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1046_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1048,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_105_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_105_final_reg_req_0;
      addr_of_105_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_105_final_reg_req_1;
      addr_of_105_final_reg_ack_1<= rack(0);
      addr_of_105_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_105_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_104_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr1_106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1073_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1073_final_reg_req_0;
      addr_of_1073_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1073_final_reg_req_1;
      addr_of_1073_final_reg_ack_1<= rack(0);
      addr_of_1073_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1073_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1072_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1099_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1099_final_reg_req_0;
      addr_of_1099_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1099_final_reg_req_1;
      addr_of_1099_final_reg_ack_1<= rack(0);
      addr_of_1099_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1099_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1098_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1100,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1125_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1125_final_reg_req_0;
      addr_of_1125_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1125_final_reg_req_1;
      addr_of_1125_final_reg_ack_1<= rack(0);
      addr_of_1125_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1125_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1124_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_112_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_112_final_reg_req_0;
      addr_of_112_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_112_final_reg_req_1;
      addr_of_112_final_reg_ack_1<= rack(0);
      addr_of_112_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_112_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_111_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr2_113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_119_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_119_final_reg_req_0;
      addr_of_119_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_119_final_reg_req_1;
      addr_of_119_final_reg_ack_1<= rack(0);
      addr_of_119_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_119_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_118_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr3_120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_126_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_126_final_reg_req_0;
      addr_of_126_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_126_final_reg_req_1;
      addr_of_126_final_reg_ack_1<= rack(0);
      addr_of_126_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_126_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_125_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr4_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1055_inst
    process(out1_681) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out1_681(15 downto 0);
      type_cast_1055_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1057_inst
    process(out2_705) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out2_705(15 downto 0);
      type_cast_1057_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1060_inst
    process(out3_729) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out3_729(15 downto 0);
      type_cast_1060_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1062_inst
    process(out4_753) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out4_753(15 downto 0);
      type_cast_1062_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1081_inst
    process(out5_777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out5_777(15 downto 0);
      type_cast_1081_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1083_inst
    process(out6_801) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out6_801(15 downto 0);
      type_cast_1083_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1086_inst
    process(out7_825) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out7_825(15 downto 0);
      type_cast_1086_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1088_inst
    process(out8_849) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out8_849(15 downto 0);
      type_cast_1088_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1107_inst
    process(out9_873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out9_873(15 downto 0);
      type_cast_1107_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1109_inst
    process(out10_897) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out10_897(15 downto 0);
      type_cast_1109_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1112_inst
    process(out11_921) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out11_921(15 downto 0);
      type_cast_1112_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1114_inst
    process(out12_945) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out12_945(15 downto 0);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1133_inst
    process(out13_969) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out13_969(15 downto 0);
      type_cast_1133_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1135_inst
    process(out14_993) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out14_993(15 downto 0);
      type_cast_1135_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1138_inst
    process(out15_1017) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out15_1017(15 downto 0);
      type_cast_1138_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1140_inst
    process(out16_1041) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out16_1041(15 downto 0);
      type_cast_1140_wire <= tmp_var; -- 
    end process;
    type_cast_1146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1146_inst_req_0;
      type_cast_1146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1146_inst_req_1;
      type_cast_1146_inst_ack_1<= rack(0);
      type_cast_1146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_404_inst
    process(sliced_v11_148) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v11_148(15 downto 0);
      a11_405 <= tmp_var; -- 
    end process;
    -- interlock type_cast_408_inst
    process(sliced_v12_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v12_152(15 downto 0);
      a12_409 <= tmp_var; -- 
    end process;
    -- interlock type_cast_412_inst
    process(sliced_v13_156) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v13_156(15 downto 0);
      a13_413 <= tmp_var; -- 
    end process;
    -- interlock type_cast_416_inst
    process(sliced_v14_160) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v14_160(15 downto 0);
      a14_417 <= tmp_var; -- 
    end process;
    -- interlock type_cast_420_inst
    process(sliced_v15_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v15_164(15 downto 0);
      a15_421 <= tmp_var; -- 
    end process;
    -- interlock type_cast_424_inst
    process(sliced_v16_168) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v16_168(15 downto 0);
      a16_425 <= tmp_var; -- 
    end process;
    -- interlock type_cast_428_inst
    process(sliced_v17_172) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v17_172(15 downto 0);
      a17_429 <= tmp_var; -- 
    end process;
    -- interlock type_cast_432_inst
    process(sliced_v18_176) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v18_176(15 downto 0);
      a18_433 <= tmp_var; -- 
    end process;
    -- interlock type_cast_436_inst
    process(sliced_v19_180) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v19_180(15 downto 0);
      a19_437 <= tmp_var; -- 
    end process;
    -- interlock type_cast_440_inst
    process(sliced_v110_184) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v110_184(15 downto 0);
      a110_441 <= tmp_var; -- 
    end process;
    -- interlock type_cast_444_inst
    process(sliced_v111_188) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v111_188(15 downto 0);
      a111_445 <= tmp_var; -- 
    end process;
    -- interlock type_cast_448_inst
    process(sliced_v112_192) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v112_192(15 downto 0);
      a112_449 <= tmp_var; -- 
    end process;
    -- interlock type_cast_452_inst
    process(sliced_v113_196) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v113_196(15 downto 0);
      a113_453 <= tmp_var; -- 
    end process;
    -- interlock type_cast_456_inst
    process(sliced_v114_200) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v114_200(15 downto 0);
      a114_457 <= tmp_var; -- 
    end process;
    -- interlock type_cast_460_inst
    process(sliced_v115_204) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v115_204(15 downto 0);
      a115_461 <= tmp_var; -- 
    end process;
    -- interlock type_cast_464_inst
    process(sliced_v116_208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v116_208(15 downto 0);
      a116_465 <= tmp_var; -- 
    end process;
    -- interlock type_cast_468_inst
    process(sliced_v21_212) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v21_212(15 downto 0);
      a21_469 <= tmp_var; -- 
    end process;
    -- interlock type_cast_472_inst
    process(sliced_v22_216) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v22_216(15 downto 0);
      a22_473 <= tmp_var; -- 
    end process;
    -- interlock type_cast_476_inst
    process(sliced_v23_220) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v23_220(15 downto 0);
      a23_477 <= tmp_var; -- 
    end process;
    -- interlock type_cast_480_inst
    process(sliced_v24_224) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v24_224(15 downto 0);
      a24_481 <= tmp_var; -- 
    end process;
    -- interlock type_cast_484_inst
    process(sliced_v25_228) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v25_228(15 downto 0);
      a25_485 <= tmp_var; -- 
    end process;
    -- interlock type_cast_488_inst
    process(sliced_v26_232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v26_232(15 downto 0);
      a26_489 <= tmp_var; -- 
    end process;
    -- interlock type_cast_492_inst
    process(sliced_v27_236) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v27_236(15 downto 0);
      a27_493 <= tmp_var; -- 
    end process;
    -- interlock type_cast_496_inst
    process(sliced_v28_240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v28_240(15 downto 0);
      a28_497 <= tmp_var; -- 
    end process;
    -- interlock type_cast_500_inst
    process(sliced_v29_244) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v29_244(15 downto 0);
      a29_501 <= tmp_var; -- 
    end process;
    -- interlock type_cast_504_inst
    process(sliced_v210_248) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v210_248(15 downto 0);
      a210_505 <= tmp_var; -- 
    end process;
    -- interlock type_cast_508_inst
    process(sliced_v211_252) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v211_252(15 downto 0);
      a211_509 <= tmp_var; -- 
    end process;
    -- interlock type_cast_512_inst
    process(sliced_v212_256) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v212_256(15 downto 0);
      a212_513 <= tmp_var; -- 
    end process;
    -- interlock type_cast_516_inst
    process(sliced_v213_260) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v213_260(15 downto 0);
      a213_517 <= tmp_var; -- 
    end process;
    -- interlock type_cast_520_inst
    process(sliced_v214_264) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v214_264(15 downto 0);
      a214_521 <= tmp_var; -- 
    end process;
    -- interlock type_cast_524_inst
    process(sliced_v215_268) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v215_268(15 downto 0);
      a215_525 <= tmp_var; -- 
    end process;
    -- interlock type_cast_528_inst
    process(sliced_v216_272) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v216_272(15 downto 0);
      a216_529 <= tmp_var; -- 
    end process;
    -- interlock type_cast_532_inst
    process(sliced_v31_276) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v31_276(15 downto 0);
      a31_533 <= tmp_var; -- 
    end process;
    -- interlock type_cast_536_inst
    process(sliced_v32_280) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v32_280(15 downto 0);
      a32_537 <= tmp_var; -- 
    end process;
    -- interlock type_cast_540_inst
    process(sliced_v33_284) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v33_284(15 downto 0);
      a33_541 <= tmp_var; -- 
    end process;
    -- interlock type_cast_544_inst
    process(sliced_v34_288) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v34_288(15 downto 0);
      a34_545 <= tmp_var; -- 
    end process;
    -- interlock type_cast_548_inst
    process(sliced_v35_292) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v35_292(15 downto 0);
      a35_549 <= tmp_var; -- 
    end process;
    -- interlock type_cast_552_inst
    process(sliced_v36_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v36_296(15 downto 0);
      a36_553 <= tmp_var; -- 
    end process;
    -- interlock type_cast_556_inst
    process(sliced_v37_300) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v37_300(15 downto 0);
      a37_557 <= tmp_var; -- 
    end process;
    -- interlock type_cast_560_inst
    process(sliced_v38_304) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v38_304(15 downto 0);
      a38_561 <= tmp_var; -- 
    end process;
    -- interlock type_cast_564_inst
    process(sliced_v39_308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v39_308(15 downto 0);
      a39_565 <= tmp_var; -- 
    end process;
    -- interlock type_cast_568_inst
    process(sliced_v310_312) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v310_312(15 downto 0);
      a310_569 <= tmp_var; -- 
    end process;
    -- interlock type_cast_572_inst
    process(sliced_v311_316) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v311_316(15 downto 0);
      a311_573 <= tmp_var; -- 
    end process;
    -- interlock type_cast_576_inst
    process(sliced_v312_320) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v312_320(15 downto 0);
      a312_577 <= tmp_var; -- 
    end process;
    -- interlock type_cast_580_inst
    process(sliced_v313_324) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v313_324(15 downto 0);
      a313_581 <= tmp_var; -- 
    end process;
    -- interlock type_cast_584_inst
    process(sliced_v314_328) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v314_328(15 downto 0);
      a314_585 <= tmp_var; -- 
    end process;
    -- interlock type_cast_588_inst
    process(sliced_v315_332) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v315_332(15 downto 0);
      a315_589 <= tmp_var; -- 
    end process;
    -- interlock type_cast_592_inst
    process(sliced_v316_336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v316_336(15 downto 0);
      a316_593 <= tmp_var; -- 
    end process;
    -- interlock type_cast_596_inst
    process(sliced_v41_340) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v41_340(15 downto 0);
      a41_597 <= tmp_var; -- 
    end process;
    -- interlock type_cast_600_inst
    process(sliced_v42_344) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v42_344(15 downto 0);
      a42_601 <= tmp_var; -- 
    end process;
    -- interlock type_cast_604_inst
    process(sliced_v43_348) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v43_348(15 downto 0);
      a43_605 <= tmp_var; -- 
    end process;
    -- interlock type_cast_608_inst
    process(sliced_v44_352) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v44_352(15 downto 0);
      a44_609 <= tmp_var; -- 
    end process;
    -- interlock type_cast_612_inst
    process(sliced_v45_356) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v45_356(15 downto 0);
      a45_613 <= tmp_var; -- 
    end process;
    -- interlock type_cast_616_inst
    process(sliced_v46_360) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v46_360(15 downto 0);
      a46_617 <= tmp_var; -- 
    end process;
    -- interlock type_cast_620_inst
    process(sliced_v47_364) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v47_364(15 downto 0);
      a47_621 <= tmp_var; -- 
    end process;
    -- interlock type_cast_624_inst
    process(sliced_v48_368) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v48_368(15 downto 0);
      a48_625 <= tmp_var; -- 
    end process;
    -- interlock type_cast_628_inst
    process(sliced_v49_372) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v49_372(15 downto 0);
      a49_629 <= tmp_var; -- 
    end process;
    -- interlock type_cast_632_inst
    process(sliced_v410_376) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v410_376(15 downto 0);
      a410_633 <= tmp_var; -- 
    end process;
    -- interlock type_cast_636_inst
    process(sliced_v411_380) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v411_380(15 downto 0);
      a411_637 <= tmp_var; -- 
    end process;
    -- interlock type_cast_640_inst
    process(sliced_v412_384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v412_384(15 downto 0);
      a412_641 <= tmp_var; -- 
    end process;
    -- interlock type_cast_644_inst
    process(sliced_v413_388) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v413_388(15 downto 0);
      a413_645 <= tmp_var; -- 
    end process;
    -- interlock type_cast_648_inst
    process(sliced_v414_392) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v414_392(15 downto 0);
      a414_649 <= tmp_var; -- 
    end process;
    -- interlock type_cast_652_inst
    process(sliced_v415_396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v415_396(15 downto 0);
      a415_653 <= tmp_var; -- 
    end process;
    -- interlock type_cast_656_inst
    process(sliced_v416_400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v416_400(15 downto 0);
      a416_657 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_1046_index_1_rename
    process(R_addr_1045_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1045_resized;
      ov(13 downto 0) := iv;
      R_addr_1045_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1046_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_1045_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1046_root_address_inst
    process(array_obj_ref_1046_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1046_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1046_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_104_index_1_rename
    process(R_addr1_103_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_103_resized;
      ov(13 downto 0) := iv;
      R_addr1_103_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_104_index_1_resize
    process(addr1_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_buffer;
      ov := iv(13 downto 0);
      R_addr1_103_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_104_root_address_inst
    process(array_obj_ref_104_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_104_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_104_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_rename
    process(ADD_u32_u32_1071_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1071_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1071_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_index_1_resize
    process(ADD_u32_u32_1071_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1071_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1071_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1072_root_address_inst
    process(array_obj_ref_1072_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1072_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1098_index_1_rename
    process(ADD_u32_u32_1097_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1097_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1097_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1098_index_1_resize
    process(ADD_u32_u32_1097_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1097_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1097_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1098_root_address_inst
    process(array_obj_ref_1098_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1098_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1098_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_111_index_1_rename
    process(R_addr2_110_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_110_resized;
      ov(13 downto 0) := iv;
      R_addr2_110_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_111_index_1_resize
    process(addr2_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_buffer;
      ov := iv(13 downto 0);
      R_addr2_110_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_111_root_address_inst
    process(array_obj_ref_111_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_111_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_111_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1124_index_1_rename
    process(ADD_u32_u32_1123_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1123_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1123_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1124_index_1_resize
    process(ADD_u32_u32_1123_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1123_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1123_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1124_root_address_inst
    process(array_obj_ref_1124_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1124_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1124_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_118_index_1_rename
    process(R_addr3_117_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_117_resized;
      ov(13 downto 0) := iv;
      R_addr3_117_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_118_index_1_resize
    process(addr3_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_buffer;
      ov := iv(13 downto 0);
      R_addr3_117_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_118_root_address_inst
    process(array_obj_ref_118_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_118_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_118_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_1_rename
    process(R_addr4_124_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr4_124_resized;
      ov(13 downto 0) := iv;
      R_addr4_124_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_index_1_resize
    process(addr4_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr4_buffer;
      ov := iv(13 downto 0);
      R_addr4_124_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_125_root_address_inst
    process(array_obj_ref_125_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_125_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_125_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1053_addr_0
    process(ptr_deref_1053_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1053_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1053_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1053_base_resize
    process(myptr5_1049_delayed_8_0_1051) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr5_1049_delayed_8_0_1051;
      ov := iv(13 downto 0);
      ptr_deref_1053_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1053_gather_scatter
    process(CONCAT_u32_u64_1064_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1064_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1053_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1053_root_address_inst
    process(ptr_deref_1053_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1053_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1053_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1079_addr_0
    process(ptr_deref_1079_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1079_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1079_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1079_base_resize
    process(myptr6_1072_delayed_8_0_1077) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr6_1072_delayed_8_0_1077;
      ov := iv(13 downto 0);
      ptr_deref_1079_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1079_gather_scatter
    process(CONCAT_u32_u64_1090_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1090_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1079_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1079_root_address_inst
    process(ptr_deref_1079_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1079_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1079_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1105_addr_0
    process(ptr_deref_1105_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1105_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1105_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1105_base_resize
    process(myptr7_1095_delayed_8_0_1103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr7_1095_delayed_8_0_1103;
      ov := iv(13 downto 0);
      ptr_deref_1105_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1105_gather_scatter
    process(CONCAT_u32_u64_1116_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1116_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1105_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1105_root_address_inst
    process(ptr_deref_1105_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1105_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1105_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1131_addr_0
    process(ptr_deref_1131_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1131_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1131_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1131_base_resize
    process(myptr8_1118_delayed_8_0_1129) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr8_1118_delayed_8_0_1129;
      ov := iv(13 downto 0);
      ptr_deref_1131_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1131_gather_scatter
    process(CONCAT_u32_u64_1142_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1142_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1131_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1131_root_address_inst
    process(ptr_deref_1131_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1131_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1131_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_addr_0
    process(ptr_deref_130_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_130_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_130_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_base_resize
    process(myptr1_106) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr1_106;
      ov := iv(13 downto 0);
      ptr_deref_130_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_gather_scatter
    process(ptr_deref_130_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_130_data_0;
      ov(255 downto 0) := iv;
      c1_131 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_root_address_inst
    process(ptr_deref_130_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_130_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_130_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_134_addr_0
    process(ptr_deref_134_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_134_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_134_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_134_base_resize
    process(myptr2_113) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr2_113;
      ov := iv(13 downto 0);
      ptr_deref_134_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_134_gather_scatter
    process(ptr_deref_134_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_134_data_0;
      ov(255 downto 0) := iv;
      c2_135 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_134_root_address_inst
    process(ptr_deref_134_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_134_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_134_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_addr_0
    process(ptr_deref_138_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_base_resize
    process(myptr3_120) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr3_120;
      ov := iv(13 downto 0);
      ptr_deref_138_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_gather_scatter
    process(ptr_deref_138_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_data_0;
      ov(255 downto 0) := iv;
      c3_139 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_root_address_inst
    process(ptr_deref_138_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_addr_0
    process(ptr_deref_142_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_142_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_base_resize
    process(myptr4_127) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr4_127;
      ov := iv(13 downto 0);
      ptr_deref_142_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_gather_scatter
    process(ptr_deref_142_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_data_0;
      ov(255 downto 0) := iv;
      c4_143 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_root_address_inst
    process(ptr_deref_142_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_142_root_address <= ov(13 downto 0);
      --
    end process;
    -- binary operator ADD_u32_u32_1071_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1070_wire_constant, tmp_var);
      ADD_u32_u32_1071_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1097_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1096_wire_constant, tmp_var);
      ADD_u32_u32_1097_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1123_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1122_wire_constant, tmp_var);
      ADD_u32_u32_1123_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1058_inst
    process(type_cast_1055_wire, type_cast_1057_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1055_wire, type_cast_1057_wire, tmp_var);
      CONCAT_u16_u32_1058_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1063_inst
    process(type_cast_1060_wire, type_cast_1062_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1060_wire, type_cast_1062_wire, tmp_var);
      CONCAT_u16_u32_1063_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1084_inst
    process(type_cast_1081_wire, type_cast_1083_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1081_wire, type_cast_1083_wire, tmp_var);
      CONCAT_u16_u32_1084_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1089_inst
    process(type_cast_1086_wire, type_cast_1088_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1086_wire, type_cast_1088_wire, tmp_var);
      CONCAT_u16_u32_1089_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1110_inst
    process(type_cast_1107_wire, type_cast_1109_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1107_wire, type_cast_1109_wire, tmp_var);
      CONCAT_u16_u32_1110_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1115_inst
    process(type_cast_1112_wire, type_cast_1114_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1112_wire, type_cast_1114_wire, tmp_var);
      CONCAT_u16_u32_1115_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1136_inst
    process(type_cast_1133_wire, type_cast_1135_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1133_wire, type_cast_1135_wire, tmp_var);
      CONCAT_u16_u32_1136_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1141_inst
    process(type_cast_1138_wire, type_cast_1140_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1138_wire, type_cast_1140_wire, tmp_var);
      CONCAT_u16_u32_1141_wire <= tmp_var; --
    end process;
    -- shared split operator group (11) : CONCAT_u32_u64_1064_inst 
    ApConcat_group_11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1058_wire & CONCAT_u16_u32_1063_wire;
      CONCAT_u32_u64_1064_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1064_inst_req_0;
      CONCAT_u32_u64_1064_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1064_inst_req_1;
      CONCAT_u32_u64_1064_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_11_gI: SplitGuardInterface generic map(name => "ApConcat_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : CONCAT_u32_u64_1090_inst 
    ApConcat_group_12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1084_wire & CONCAT_u16_u32_1089_wire;
      CONCAT_u32_u64_1090_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1090_inst_req_0;
      CONCAT_u32_u64_1090_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1090_inst_req_1;
      CONCAT_u32_u64_1090_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_12_gI: SplitGuardInterface generic map(name => "ApConcat_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : CONCAT_u32_u64_1116_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1110_wire & CONCAT_u16_u32_1115_wire;
      CONCAT_u32_u64_1116_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1116_inst_req_0;
      CONCAT_u32_u64_1116_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1116_inst_req_1;
      CONCAT_u32_u64_1116_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_1142_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1136_wire & CONCAT_u16_u32_1141_wire;
      CONCAT_u32_u64_1142_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1142_inst_req_0;
      CONCAT_u32_u64_1142_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1142_inst_req_1;
      CONCAT_u32_u64_1142_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator SGT_i16_u1_1005_inst
    process(a315_589, a415_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a315_589, a415_653, tmp_var);
      SGT_i16_u1_1005_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1013_inst
    process(t151_1001, t152_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t151_1001, t152_1009, tmp_var);
      SGT_i16_u1_1013_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1021_inst
    process(a116_465, a216_529) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a116_465, a216_529, tmp_var);
      SGT_i16_u1_1021_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1029_inst
    process(a316_593, a416_657) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a316_593, a416_657, tmp_var);
      SGT_i16_u1_1029_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1037_inst
    process(t161_1025, t162_1033) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t161_1025, t162_1033, tmp_var);
      SGT_i16_u1_1037_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_661_inst
    process(a11_405, a21_469) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_405, a21_469, tmp_var);
      SGT_i16_u1_661_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_669_inst
    process(a31_533, a41_597) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_533, a41_597, tmp_var);
      SGT_i16_u1_669_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_677_inst
    process(t11_665, t12_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_665, t12_673, tmp_var);
      SGT_i16_u1_677_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_685_inst
    process(a12_409, a22_473) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_409, a22_473, tmp_var);
      SGT_i16_u1_685_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_693_inst
    process(a32_537, a42_601) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_537, a42_601, tmp_var);
      SGT_i16_u1_693_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_701_inst
    process(t21_689, t22_697) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_689, t22_697, tmp_var);
      SGT_i16_u1_701_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_709_inst
    process(a13_413, a23_477) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_413, a23_477, tmp_var);
      SGT_i16_u1_709_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_717_inst
    process(a33_541, a43_605) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_541, a43_605, tmp_var);
      SGT_i16_u1_717_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_725_inst
    process(t31_713, t32_721) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_713, t32_721, tmp_var);
      SGT_i16_u1_725_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_733_inst
    process(a14_417, a24_481) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_417, a24_481, tmp_var);
      SGT_i16_u1_733_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_741_inst
    process(a34_545, a44_609) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_545, a44_609, tmp_var);
      SGT_i16_u1_741_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_749_inst
    process(t41_737, t42_745) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_737, t42_745, tmp_var);
      SGT_i16_u1_749_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_757_inst
    process(a15_421, a25_485) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a15_421, a25_485, tmp_var);
      SGT_i16_u1_757_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_765_inst
    process(a35_549, a45_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a35_549, a45_613, tmp_var);
      SGT_i16_u1_765_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_773_inst
    process(t51_761, t52_769) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t51_761, t52_769, tmp_var);
      SGT_i16_u1_773_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_781_inst
    process(a16_425, a26_489) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a16_425, a26_489, tmp_var);
      SGT_i16_u1_781_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_789_inst
    process(a36_553, a46_617) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a36_553, a46_617, tmp_var);
      SGT_i16_u1_789_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_797_inst
    process(t61_785, t62_793) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t61_785, t62_793, tmp_var);
      SGT_i16_u1_797_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_805_inst
    process(a17_429, a27_493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a17_429, a27_493, tmp_var);
      SGT_i16_u1_805_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_813_inst
    process(a37_557, a47_621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a37_557, a47_621, tmp_var);
      SGT_i16_u1_813_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_821_inst
    process(t71_809, t72_817) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t71_809, t72_817, tmp_var);
      SGT_i16_u1_821_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_829_inst
    process(a18_433, a28_497) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a18_433, a28_497, tmp_var);
      SGT_i16_u1_829_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_837_inst
    process(a38_561, a48_625) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a38_561, a48_625, tmp_var);
      SGT_i16_u1_837_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_845_inst
    process(t81_833, t82_841) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t81_833, t82_841, tmp_var);
      SGT_i16_u1_845_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_853_inst
    process(a19_437, a29_501) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a19_437, a29_501, tmp_var);
      SGT_i16_u1_853_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_861_inst
    process(a39_565, a49_629) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a39_565, a49_629, tmp_var);
      SGT_i16_u1_861_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_869_inst
    process(t91_857, t92_865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t91_857, t92_865, tmp_var);
      SGT_i16_u1_869_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_877_inst
    process(a110_441, a210_505) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a110_441, a210_505, tmp_var);
      SGT_i16_u1_877_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_885_inst
    process(a310_569, a410_633) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a310_569, a410_633, tmp_var);
      SGT_i16_u1_885_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_893_inst
    process(t101_881, t102_889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t101_881, t102_889, tmp_var);
      SGT_i16_u1_893_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_901_inst
    process(a111_445, a211_509) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a111_445, a211_509, tmp_var);
      SGT_i16_u1_901_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_909_inst
    process(a311_573, a411_637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a311_573, a411_637, tmp_var);
      SGT_i16_u1_909_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_917_inst
    process(t111_905, t112_913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t111_905, t112_913, tmp_var);
      SGT_i16_u1_917_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_925_inst
    process(a112_449, a212_513) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a112_449, a212_513, tmp_var);
      SGT_i16_u1_925_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_933_inst
    process(a312_577, a412_641) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a312_577, a412_641, tmp_var);
      SGT_i16_u1_933_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_941_inst
    process(t121_929, t122_937) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t121_929, t122_937, tmp_var);
      SGT_i16_u1_941_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_949_inst
    process(a113_453, a213_517) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a113_453, a213_517, tmp_var);
      SGT_i16_u1_949_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_957_inst
    process(a313_581, a413_645) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a313_581, a413_645, tmp_var);
      SGT_i16_u1_957_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_965_inst
    process(t131_953, t132_961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t131_953, t132_961, tmp_var);
      SGT_i16_u1_965_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_973_inst
    process(a114_457, a214_521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a114_457, a214_521, tmp_var);
      SGT_i16_u1_973_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_981_inst
    process(a314_585, a414_649) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a314_585, a414_649, tmp_var);
      SGT_i16_u1_981_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_989_inst
    process(t141_977, t142_985) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t141_977, t142_985, tmp_var);
      SGT_i16_u1_989_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_997_inst
    process(a115_461, a215_525) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a115_461, a215_525, tmp_var);
      SGT_i16_u1_997_wire <= tmp_var; --
    end process;
    -- shared split operator group (63) : array_obj_ref_1046_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_1045_scaled;
      array_obj_ref_1046_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1046_index_offset_req_0;
      array_obj_ref_1046_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1046_index_offset_req_1;
      array_obj_ref_1046_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : array_obj_ref_104_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr1_103_scaled;
      array_obj_ref_104_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_104_index_offset_req_0;
      array_obj_ref_104_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_104_index_offset_req_1;
      array_obj_ref_104_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : array_obj_ref_1072_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1071_scaled;
      array_obj_ref_1072_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1072_index_offset_req_0;
      array_obj_ref_1072_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1072_index_offset_req_1;
      array_obj_ref_1072_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_1098_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1097_scaled;
      array_obj_ref_1098_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1098_index_offset_req_0;
      array_obj_ref_1098_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1098_index_offset_req_1;
      array_obj_ref_1098_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : array_obj_ref_111_index_offset 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr2_110_scaled;
      array_obj_ref_111_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_111_index_offset_req_0;
      array_obj_ref_111_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_111_index_offset_req_1;
      array_obj_ref_111_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_67_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : array_obj_ref_1124_index_offset 
    ApIntAdd_group_68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1123_scaled;
      array_obj_ref_1124_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1124_index_offset_req_0;
      array_obj_ref_1124_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1124_index_offset_req_1;
      array_obj_ref_1124_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_68_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_68_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : array_obj_ref_118_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr3_117_scaled;
      array_obj_ref_118_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_118_index_offset_req_0;
      array_obj_ref_118_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_118_index_offset_req_1;
      array_obj_ref_118_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_125_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr4_124_scaled;
      array_obj_ref_125_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_125_index_offset_req_0;
      array_obj_ref_125_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_125_index_offset_req_1;
      array_obj_ref_125_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared load operator group (0) : ptr_deref_130_load_0 ptr_deref_134_load_0 ptr_deref_138_load_0 ptr_deref_142_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_130_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_134_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_138_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_142_load_0_req_0;
      ptr_deref_130_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_134_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_138_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_142_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_130_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_134_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_138_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_142_load_0_req_1;
      ptr_deref_130_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_134_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_138_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_142_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_130_word_address_0 & ptr_deref_134_word_address_0 & ptr_deref_138_word_address_0 & ptr_deref_142_word_address_0;
      ptr_deref_130_data_0 <= data_out(1023 downto 768);
      ptr_deref_134_data_0 <= data_out(767 downto 512);
      ptr_deref_138_data_0 <= data_out(511 downto 256);
      ptr_deref_142_data_0 <= data_out(255 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 256,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(255 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1053_store_0 ptr_deref_1079_store_0 ptr_deref_1105_store_0 ptr_deref_1131_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 15, 2 => 15, 1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_1053_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1079_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1105_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1131_store_0_req_0;
      ptr_deref_1053_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1079_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1105_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1131_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_1053_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1079_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1105_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1131_store_0_req_1;
      ptr_deref_1053_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1079_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1105_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1131_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1053_word_address_0 & ptr_deref_1079_word_address_0 & ptr_deref_1105_word_address_0 & ptr_deref_1131_word_address_0;
      data_in <= ptr_deref_1053_data_0 & ptr_deref_1079_data_0 & ptr_deref_1105_data_0 & ptr_deref_1131_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2178_start: Boolean;
  signal sendB_CP_2178_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_1214_index_offset_req_1 : boolean;
  signal array_obj_ref_1214_index_offset_ack_1 : boolean;
  signal type_cast_1185_inst_req_0 : boolean;
  signal if_stmt_1158_branch_req_0 : boolean;
  signal type_cast_1185_inst_ack_0 : boolean;
  signal if_stmt_1158_branch_ack_0 : boolean;
  signal type_cast_1185_inst_ack_1 : boolean;
  signal if_stmt_1158_branch_ack_1 : boolean;
  signal array_obj_ref_1214_index_offset_req_0 : boolean;
  signal array_obj_ref_1214_index_offset_ack_0 : boolean;
  signal type_cast_1185_inst_req_1 : boolean;
  signal ptr_deref_1219_load_0_req_0 : boolean;
  signal ptr_deref_1219_load_0_ack_0 : boolean;
  signal addr_of_1215_final_reg_req_1 : boolean;
  signal ptr_deref_1219_load_0_req_1 : boolean;
  signal ptr_deref_1219_load_0_ack_1 : boolean;
  signal addr_of_1215_final_reg_req_0 : boolean;
  signal addr_of_1215_final_reg_ack_0 : boolean;
  signal addr_of_1215_final_reg_ack_1 : boolean;
  signal type_cast_1265_inst_req_0 : boolean;
  signal type_cast_1265_inst_ack_0 : boolean;
  signal type_cast_1265_inst_req_1 : boolean;
  signal type_cast_1265_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1267_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1267_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1267_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1267_inst_ack_1 : boolean;
  signal type_cast_1272_inst_req_0 : boolean;
  signal type_cast_1272_inst_ack_0 : boolean;
  signal type_cast_1272_inst_req_1 : boolean;
  signal type_cast_1272_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1274_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1274_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1274_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1274_inst_ack_1 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1281_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1281_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1281_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1281_inst_ack_1 : boolean;
  signal type_cast_1286_inst_req_0 : boolean;
  signal type_cast_1286_inst_ack_0 : boolean;
  signal type_cast_1286_inst_req_1 : boolean;
  signal type_cast_1286_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1288_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1288_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1288_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1288_inst_ack_1 : boolean;
  signal type_cast_1293_inst_req_0 : boolean;
  signal type_cast_1293_inst_ack_0 : boolean;
  signal type_cast_1293_inst_req_1 : boolean;
  signal type_cast_1293_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1295_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1295_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1295_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1295_inst_ack_1 : boolean;
  signal type_cast_1300_inst_req_0 : boolean;
  signal type_cast_1300_inst_ack_0 : boolean;
  signal type_cast_1300_inst_req_1 : boolean;
  signal type_cast_1300_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1302_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1302_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1302_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1302_inst_ack_1 : boolean;
  signal type_cast_1307_inst_req_0 : boolean;
  signal type_cast_1307_inst_ack_0 : boolean;
  signal type_cast_1307_inst_req_1 : boolean;
  signal type_cast_1307_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1309_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1309_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1309_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1309_inst_ack_1 : boolean;
  signal type_cast_1314_inst_req_0 : boolean;
  signal type_cast_1314_inst_ack_0 : boolean;
  signal type_cast_1314_inst_req_1 : boolean;
  signal type_cast_1314_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1316_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1316_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1316_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1316_inst_ack_1 : boolean;
  signal if_stmt_1330_branch_req_0 : boolean;
  signal if_stmt_1330_branch_ack_1 : boolean;
  signal if_stmt_1330_branch_ack_0 : boolean;
  signal phi_stmt_1202_req_0 : boolean;
  signal type_cast_1208_inst_req_0 : boolean;
  signal type_cast_1208_inst_ack_0 : boolean;
  signal type_cast_1208_inst_req_1 : boolean;
  signal type_cast_1208_inst_ack_1 : boolean;
  signal phi_stmt_1202_req_1 : boolean;
  signal phi_stmt_1202_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2178_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2178_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2178_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2178_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2178: Block -- control-path 
    signal sendB_CP_2178_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendB_CP_2178_elements(0) <= sendB_CP_2178_start;
    sendB_CP_2178_symbol <= sendB_CP_2178_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/assign_stmt_1157/$exit
      -- CP-element group 0: 	 branch_block_stmt_1151/assign_stmt_1157__exit__
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1151/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/assign_stmt_1157/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1151/if_stmt_1158_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_1151/assign_stmt_1157__entry__
      -- CP-element group 0: 	 branch_block_stmt_1151/R_cmp76_1159_place
      -- CP-element group 0: 	 branch_block_stmt_1151/branch_block_stmt_1151__entry__
      -- 
    branch_req_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(0), ack => if_stmt_1158_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/$entry
      -- CP-element group 1: 	 branch_block_stmt_1151/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1151/merge_stmt_1164__exit__
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199__entry__
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_1151/if_stmt_1158_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_1151/if_stmt_1158_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1151/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1151/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_1151/merge_stmt_1164_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_1151/merge_stmt_1164_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_1151/merge_stmt_1164_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_1151/merge_stmt_1164_PhiAck/dummy
      -- 
    if_choice_transition_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1158_branch_ack_1, ack => sendB_CP_2178_elements(1)); -- 
    rr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(1), ack => type_cast_1185_inst_req_0); -- 
    cr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(1), ack => type_cast_1185_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1151/if_stmt_1158_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1151/if_stmt_1158_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1151/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_1151/entry_forx_xend_PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_1151/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1158_branch_ack_0, ack => sendB_CP_2178_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Sample/$exit
      -- 
    ra_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1185_inst_ack_0, ack => sendB_CP_2178_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/$exit
      -- CP-element group 4: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199__exit__
      -- CP-element group 4: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_1151/assign_stmt_1170_to_assign_stmt_1199/type_cast_1185_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/$entry
      -- CP-element group 4: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/$entry
      -- 
    ca_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1185_inst_ack_1, ack => sendB_CP_2178_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Sample/ack
      -- 
    ack_2273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1214_index_offset_ack_0, ack => sendB_CP_2178_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_request/req
      -- CP-element group 6: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_request/$entry
      -- 
    ack_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1214_index_offset_ack_1, ack => sendB_CP_2178_elements(6)); -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(6), ack => addr_of_1215_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_request/ack
      -- CP-element group 7: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_request/$exit
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1215_final_reg_ack_0, ack => sendB_CP_2178_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/word_0/rr
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_sample_start_
      -- 
    ack_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1215_final_reg_ack_1, ack => sendB_CP_2178_elements(8)); -- 
    rr_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(8), ack => ptr_deref_1219_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_sample_completed_
      -- 
    ra_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1219_load_0_ack_0, ack => sendB_CP_2178_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	30 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/ptr_deref_1219_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/ptr_deref_1219_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/ptr_deref_1219_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/ptr_deref_1219_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Sample/rr
      -- 
    ca_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1219_load_0_ack_1, ack => sendB_CP_2178_elements(10)); -- 
    rr_2351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1265_inst_req_0); -- 
    rr_2379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1272_inst_req_0); -- 
    rr_2407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1279_inst_req_0); -- 
    rr_2435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1286_inst_req_0); -- 
    rr_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1293_inst_req_0); -- 
    rr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1300_inst_req_0); -- 
    rr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1307_inst_req_0); -- 
    rr_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(10), ack => type_cast_1314_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Sample/ra
      -- 
    ra_2352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_0, ack => sendB_CP_2178_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Sample/req
      -- 
    ca_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1265_inst_ack_1, ack => sendB_CP_2178_elements(12)); -- 
    req_2365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(12), ack => WPIPE_maxpool_output_pipe_1267_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Update/req
      -- 
    ack_2366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1267_inst_ack_0, ack => sendB_CP_2178_elements(13)); -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(13), ack => WPIPE_maxpool_output_pipe_1267_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1267_Update/ack
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1267_inst_ack_1, ack => sendB_CP_2178_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Sample/ra
      -- 
    ra_2380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_0, ack => sendB_CP_2178_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Update/ca
      -- 
    ca_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1272_inst_ack_1, ack => sendB_CP_2178_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Sample/req
      -- 
    req_2393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(17), ack => WPIPE_maxpool_output_pipe_1274_inst_req_0); -- 
    sendB_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(14) & sendB_CP_2178_elements(16);
      gj_sendB_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Update/req
      -- 
    ack_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1274_inst_ack_0, ack => sendB_CP_2178_elements(18)); -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(18), ack => WPIPE_maxpool_output_pipe_1274_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1274_Update/ack
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1274_inst_ack_1, ack => sendB_CP_2178_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Sample/ra
      -- 
    ra_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => sendB_CP_2178_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	58 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Update/ca
      -- 
    ca_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => sendB_CP_2178_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Sample/req
      -- 
    req_2421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(22), ack => WPIPE_maxpool_output_pipe_1281_inst_req_0); -- 
    sendB_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(19) & sendB_CP_2178_elements(21);
      gj_sendB_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Sample/ack
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Update/req
      -- 
    ack_2422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1281_inst_ack_0, ack => sendB_CP_2178_elements(23)); -- 
    req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(23), ack => WPIPE_maxpool_output_pipe_1281_inst_req_1); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1281_Update/ack
      -- 
    ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1281_inst_ack_1, ack => sendB_CP_2178_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Sample/ra
      -- 
    ra_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_0, ack => sendB_CP_2178_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Update/ca
      -- 
    ca_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1286_inst_ack_1, ack => sendB_CP_2178_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Sample/req
      -- 
    req_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(27), ack => WPIPE_maxpool_output_pipe_1288_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(24) & sendB_CP_2178_elements(26);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Update/req
      -- 
    ack_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1288_inst_ack_0, ack => sendB_CP_2178_elements(28)); -- 
    req_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(28), ack => WPIPE_maxpool_output_pipe_1288_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1288_Update/ack
      -- 
    ack_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1288_inst_ack_1, ack => sendB_CP_2178_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Sample/ra
      -- 
    ra_2464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1293_inst_ack_0, ack => sendB_CP_2178_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	58 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Update/ca
      -- 
    ca_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1293_inst_ack_1, ack => sendB_CP_2178_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Sample/req
      -- 
    req_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(32), ack => WPIPE_maxpool_output_pipe_1295_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(29) & sendB_CP_2178_elements(31);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Update/req
      -- 
    ack_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1295_inst_ack_0, ack => sendB_CP_2178_elements(33)); -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(33), ack => WPIPE_maxpool_output_pipe_1295_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1295_Update/ack
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1295_inst_ack_1, ack => sendB_CP_2178_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Sample/ra
      -- 
    ra_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_0, ack => sendB_CP_2178_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	58 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Update/ca
      -- 
    ca_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1300_inst_ack_1, ack => sendB_CP_2178_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Sample/req
      -- 
    req_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(37), ack => WPIPE_maxpool_output_pipe_1302_inst_req_0); -- 
    sendB_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(34) & sendB_CP_2178_elements(36);
      gj_sendB_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Update/req
      -- 
    ack_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1302_inst_ack_0, ack => sendB_CP_2178_elements(38)); -- 
    req_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(38), ack => WPIPE_maxpool_output_pipe_1302_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1302_Update/ack
      -- 
    ack_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1302_inst_ack_1, ack => sendB_CP_2178_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Sample/ra
      -- 
    ra_2520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1307_inst_ack_0, ack => sendB_CP_2178_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Update/ca
      -- 
    ca_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1307_inst_ack_1, ack => sendB_CP_2178_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Sample/req
      -- 
    req_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(42), ack => WPIPE_maxpool_output_pipe_1309_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(39) & sendB_CP_2178_elements(41);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Update/req
      -- 
    ack_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1309_inst_ack_0, ack => sendB_CP_2178_elements(43)); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(43), ack => WPIPE_maxpool_output_pipe_1309_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1309_Update/ack
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1309_inst_ack_1, ack => sendB_CP_2178_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Sample/ra
      -- 
    ra_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1314_inst_ack_0, ack => sendB_CP_2178_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	58 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Update/ca
      -- 
    ca_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1314_inst_ack_1, ack => sendB_CP_2178_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Sample/req
      -- 
    req_2561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(47), ack => WPIPE_maxpool_output_pipe_1316_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(44) & sendB_CP_2178_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Update/req
      -- 
    ack_2562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1316_inst_ack_0, ack => sendB_CP_2178_elements(48)); -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(48), ack => WPIPE_maxpool_output_pipe_1316_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/WPIPE_maxpool_output_pipe_1316_Update/ack
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1316_inst_ack_1, ack => sendB_CP_2178_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329__exit__
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330__entry__
      -- CP-element group 50: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/$exit
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_1151/R_exitcond1_1331_place
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1151/if_stmt_1330_else_link/$entry
      -- 
    branch_req_2575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(50), ack => if_stmt_1330_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(5) & sendB_CP_2178_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_1151/merge_stmt_1336__exit__
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1151/merge_stmt_1336_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_1151/merge_stmt_1336_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_1151/if_stmt_1330_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1151/if_stmt_1330_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1151/merge_stmt_1336_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1151/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1151/merge_stmt_1336_PhiReqMerge
      -- 
    if_choice_transition_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1330_branch_ack_1, ack => sendB_CP_2178_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_1151/if_stmt_1330_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1151/if_stmt_1330_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1330_branch_ack_0, ack => sendB_CP_2178_elements(52)); -- 
    rr_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(52), ack => type_cast_1208_inst_req_0); -- 
    cr_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(52), ack => type_cast_1208_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/$exit
      -- CP-element group 53: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1206_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_1151/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_req
      -- 
    phi_stmt_1202_req_2609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1202_req_2609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(53), ack => phi_stmt_1202_req_0); -- 
    -- Element group sendB_CP_2178_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendB_CP_2178_elements(4), ack => sendB_CP_2178_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Sample/ra
      -- 
    ra_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_0, ack => sendB_CP_2178_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/Update/ca
      -- 
    ca_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_1, ack => sendB_CP_2178_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/$exit
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/$exit
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_sources/type_cast_1208/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_1151/forx_xbody_forx_xbody_PhiReq/phi_stmt_1202/phi_stmt_1202_req
      -- 
    phi_stmt_1202_req_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1202_req_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(56), ack => phi_stmt_1202_req_1); -- 
    sendB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2178_elements(54) & sendB_CP_2178_elements(55);
      gj_sendB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2178_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1151/merge_stmt_1201_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1151/merge_stmt_1201_PhiAck/$entry
      -- 
    sendB_CP_2178_elements(57) <= OrReduce(sendB_CP_2178_elements(53) & sendB_CP_2178_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	21 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	31 
    -- CP-element group 58: 	36 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	46 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_1151/merge_stmt_1201__exit__
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329__entry__
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/addr_of_1215_complete/req
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/ptr_deref_1219_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/array_obj_ref_1214_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1265_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1272_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1279_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1286_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1293_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1300_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1307_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1151/assign_stmt_1216_to_assign_stmt_1329/type_cast_1314_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1151/merge_stmt_1201_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1151/merge_stmt_1201_PhiAck/phi_stmt_1202_ack
      -- 
    phi_stmt_1202_ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1202_ack_0, ack => sendB_CP_2178_elements(58)); -- 
    req_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => array_obj_ref_1214_index_offset_req_1); -- 
    req_2272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => array_obj_ref_1214_index_offset_req_0); -- 
    req_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => addr_of_1215_final_reg_req_1); -- 
    cr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => ptr_deref_1219_load_0_req_1); -- 
    cr_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1265_inst_req_1); -- 
    cr_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1272_inst_req_1); -- 
    cr_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1279_inst_req_1); -- 
    cr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1286_inst_req_1); -- 
    cr_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1293_inst_req_1); -- 
    cr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1300_inst_req_1); -- 
    cr_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1307_inst_req_1); -- 
    cr_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2178_elements(58), ack => type_cast_1314_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1340__exit__
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1340_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1340_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1151/return__
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_1151/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1151/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1151/branch_block_stmt_1151__exit__
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1340_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1151/$exit
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1338__exit__
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1338_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1340_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1338_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1338_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1151/merge_stmt_1338_PhiReqMerge
      -- 
    sendB_CP_2178_elements(59) <= OrReduce(sendB_CP_2178_elements(2) & sendB_CP_2178_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1213_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1213_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1214_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1216 : std_logic_vector(31 downto 0);
    signal cmp76_1157 : std_logic_vector(0 downto 0);
    signal conv52_1266 : std_logic_vector(7 downto 0);
    signal conv55_1273 : std_logic_vector(7 downto 0);
    signal conv58_1280 : std_logic_vector(7 downto 0);
    signal conv61_1287 : std_logic_vector(7 downto 0);
    signal conv64_1294 : std_logic_vector(7 downto 0);
    signal conv67_1301 : std_logic_vector(7 downto 0);
    signal conv70_1308 : std_logic_vector(7 downto 0);
    signal conv73_1315 : std_logic_vector(7 downto 0);
    signal exitcond1_1329 : std_logic_vector(0 downto 0);
    signal iNsTr_1_1186 : std_logic_vector(63 downto 0);
    signal indvar_1202 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1324 : std_logic_vector(63 downto 0);
    signal ptr_deref_1219_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1219_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1219_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_1232 : std_logic_vector(63 downto 0);
    signal shr21_1238 : std_logic_vector(63 downto 0);
    signal shr27_1244 : std_logic_vector(63 downto 0);
    signal shr33_1250 : std_logic_vector(63 downto 0);
    signal shr39_1256 : std_logic_vector(63 downto 0);
    signal shr45_1262 : std_logic_vector(63 downto 0);
    signal shr9_1226 : std_logic_vector(63 downto 0);
    signal shr_1170 : std_logic_vector(31 downto 0);
    signal shrx_xop_1182 : std_logic_vector(31 downto 0);
    signal tmp4_1220 : std_logic_vector(63 downto 0);
    signal tmp80_1199 : std_logic_vector(63 downto 0);
    signal tmp_1176 : std_logic_vector(0 downto 0);
    signal type_cast_1155_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1174_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1190_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1208_wire : std_logic_vector(63 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1230_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1242_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1248_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1254_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1192 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1214_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1214_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1214_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1214_resized_base_address <= "00000000000000";
    ptr_deref_1219_word_offset_0 <= "00000000000000";
    type_cast_1155_wire_constant <= "00000000000000000000000000000011";
    type_cast_1168_wire_constant <= "00000000000000000000000000000010";
    type_cast_1174_wire_constant <= "00000000000000000000000000000001";
    type_cast_1180_wire_constant <= "11111111111111111111111111111111";
    type_cast_1190_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1230_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1242_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1248_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1260_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1322_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1202: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1206_wire_constant & type_cast_1208_wire;
      req <= phi_stmt_1202_req_0 & phi_stmt_1202_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1202",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1202_ack_0,
          idata => idata,
          odata => indvar_1202,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1202
    -- flow-through select operator MUX_1198_inst
    tmp80_1199 <= xx_xop_1192 when (tmp_1176(0) /=  '0') else type_cast_1197_wire_constant;
    addr_of_1215_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1215_final_reg_req_0;
      addr_of_1215_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1215_final_reg_req_1;
      addr_of_1215_final_reg_ack_1<= rack(0);
      addr_of_1215_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1215_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1214_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1185_inst_req_0;
      type_cast_1185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1185_inst_req_1;
      type_cast_1185_inst_ack_1<= rack(0);
      type_cast_1185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_1182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_1186,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1208_inst_req_0;
      type_cast_1208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1208_inst_req_1;
      type_cast_1208_inst_ack_1<= rack(0);
      type_cast_1208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1208_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1265_inst_req_0;
      type_cast_1265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1265_inst_req_1;
      type_cast_1265_inst_ack_1<= rack(0);
      type_cast_1265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1272_inst_req_0;
      type_cast_1272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1272_inst_req_1;
      type_cast_1272_inst_ack_1<= rack(0);
      type_cast_1272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_1273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1286_inst_req_0;
      type_cast_1286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1286_inst_req_1;
      type_cast_1286_inst_ack_1<= rack(0);
      type_cast_1286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_1244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1293_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1293_inst_req_0;
      type_cast_1293_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1293_inst_req_1;
      type_cast_1293_inst_ack_1<= rack(0);
      type_cast_1293_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1293_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_1238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1294,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1300_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1300_inst_req_0;
      type_cast_1300_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1300_inst_req_1;
      type_cast_1300_inst_ack_1<= rack(0);
      type_cast_1300_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1300_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_1301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1307_inst_req_0;
      type_cast_1307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1307_inst_req_1;
      type_cast_1307_inst_ack_1<= rack(0);
      type_cast_1307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_1226,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1314_inst_req_0;
      type_cast_1314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1314_inst_req_1;
      type_cast_1314_inst_ack_1<= rack(0);
      type_cast_1314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_1220,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1214_index_1_rename
    process(R_indvar_1213_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1213_resized;
      ov(13 downto 0) := iv;
      R_indvar_1213_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1214_index_1_resize
    process(indvar_1202) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1202;
      ov := iv(13 downto 0);
      R_indvar_1213_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1214_root_address_inst
    process(array_obj_ref_1214_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1214_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1214_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_addr_0
    process(ptr_deref_1219_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1219_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1219_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_base_resize
    process(arrayidx_1216) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1216;
      ov := iv(13 downto 0);
      ptr_deref_1219_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_gather_scatter
    process(ptr_deref_1219_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1219_data_0;
      ov(63 downto 0) := iv;
      tmp4_1220 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1219_root_address_inst
    process(ptr_deref_1219_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1219_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1219_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1158_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp76_1157;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1158_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1158_branch_req_0,
          ack0 => if_stmt_1158_branch_ack_0,
          ack1 => if_stmt_1158_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1330_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1329;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1330_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1330_branch_req_0,
          ack0 => if_stmt_1330_branch_ack_0,
          ack1 => if_stmt_1330_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1181_inst
    process(shr_1170) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_1170, type_cast_1180_wire_constant, tmp_var);
      shrx_xop_1182 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1191_inst
    process(iNsTr_1_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_1186, type_cast_1190_wire_constant, tmp_var);
      xx_xop_1192 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1323_inst
    process(indvar_1202) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1202, type_cast_1322_wire_constant, tmp_var);
      indvarx_xnext_1324 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1328_inst
    process(indvarx_xnext_1324, tmp80_1199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1324, tmp80_1199, tmp_var);
      exitcond1_1329 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1169_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_1168_wire_constant, tmp_var);
      shr_1170 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1225_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1224_wire_constant, tmp_var);
      shr9_1226 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1231_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1230_wire_constant, tmp_var);
      shr15_1232 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1237_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1236_wire_constant, tmp_var);
      shr21_1238 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1243_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1242_wire_constant, tmp_var);
      shr27_1244 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1249_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1248_wire_constant, tmp_var);
      shr33_1250 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1255_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1254_wire_constant, tmp_var);
      shr39_1256 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1261_inst
    process(tmp4_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1220, type_cast_1260_wire_constant, tmp_var);
      shr45_1262 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1156_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_1155_wire_constant, tmp_var);
      cmp76_1157 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1175_inst
    process(shr_1170) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1170, type_cast_1174_wire_constant, tmp_var);
      tmp_1176 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_1214_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1213_scaled;
      array_obj_ref_1214_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1214_index_offset_req_0;
      array_obj_ref_1214_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1214_index_offset_req_1;
      array_obj_ref_1214_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_1219_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1219_load_0_req_0;
      ptr_deref_1219_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1219_load_0_req_1;
      ptr_deref_1219_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1219_word_address_0;
      ptr_deref_1219_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1274_inst WPIPE_maxpool_output_pipe_1302_inst WPIPE_maxpool_output_pipe_1316_inst WPIPE_maxpool_output_pipe_1295_inst WPIPE_maxpool_output_pipe_1309_inst WPIPE_maxpool_output_pipe_1288_inst WPIPE_maxpool_output_pipe_1281_inst WPIPE_maxpool_output_pipe_1267_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1274_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1302_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1316_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1295_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1309_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1288_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1281_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1267_inst_req_0;
      WPIPE_maxpool_output_pipe_1274_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1302_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1316_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1295_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1309_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1288_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1281_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1267_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1274_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1302_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1316_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1295_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1309_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1288_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1281_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1267_inst_req_1;
      WPIPE_maxpool_output_pipe_1274_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1302_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1316_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1295_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1309_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1288_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1281_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1267_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv55_1273 & conv67_1301 & conv73_1315 & conv64_1294 & conv70_1308 & conv61_1287 & conv58_1280 & conv52_1266;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_321_start: Boolean;
  signal timer_CP_321_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_90_load_0_req_0 : boolean;
  signal LOAD_count_90_load_0_ack_0 : boolean;
  signal LOAD_count_90_load_0_req_1 : boolean;
  signal LOAD_count_90_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_321_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_321_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_321_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_321_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_321: Block -- control-path 
    signal timer_CP_321_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_321_elements(0) <= timer_CP_321_start;
    timer_CP_321_symbol <= timer_CP_321_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_91/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_sample_start_
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_update_start_
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Update/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/word_0/cr
      -- 
    cr_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_321_elements(0), ack => LOAD_count_90_load_0_req_1); -- 
    rr_342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_321_elements(0), ack => LOAD_count_90_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_91/LOAD_count_90_sample_completed_
      -- CP-element group 1: 	 assign_stmt_91/LOAD_count_90_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_91/LOAD_count_90_Sample/word_access_start/word_0/ra
      -- 
    ra_343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_90_load_0_ack_0, ack => timer_CP_321_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_91/$exit
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_update_completed_
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/$exit
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/LOAD_count_90_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/LOAD_count_90_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/LOAD_count_90_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_91/LOAD_count_90_Update/LOAD_count_90_Merge/merge_ack
      -- 
    ca_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_90_load_0_ack_1, ack => timer_CP_321_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_90_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_90_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_90_word_address_0 <= "0";
    -- equivalence LOAD_count_90_gather_scatter
    process(LOAD_count_90_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_90_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_90_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_90_load_0_req_0;
      LOAD_count_90_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_90_load_0_req_1;
      LOAD_count_90_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_90_word_address_0;
      LOAD_count_90_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3718_start: Boolean;
  signal timerDaemon_CP_3718_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1874_branch_req_0 : boolean;
  signal phi_stmt_1876_req_1 : boolean;
  signal phi_stmt_1876_req_0 : boolean;
  signal phi_stmt_1876_ack_0 : boolean;
  signal ADD_u64_u64_1882_inst_req_0 : boolean;
  signal ADD_u64_u64_1882_inst_ack_0 : boolean;
  signal ADD_u64_u64_1882_inst_req_1 : boolean;
  signal ADD_u64_u64_1882_inst_ack_1 : boolean;
  signal STORE_count_1884_store_0_req_0 : boolean;
  signal STORE_count_1884_store_0_ack_0 : boolean;
  signal STORE_count_1884_store_0_req_1 : boolean;
  signal STORE_count_1884_store_0_ack_1 : boolean;
  signal do_while_stmt_1874_branch_ack_0 : boolean;
  signal do_while_stmt_1874_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3718_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3718_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3718_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3718_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3718: Block -- control-path 
    signal timerDaemon_CP_3718_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3718_elements(0) <= timerDaemon_CP_3718_start;
    timerDaemon_CP_3718_symbol <= timerDaemon_CP_3718_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1873/$entry
      -- CP-element group 0: 	 branch_block_stmt_1873/branch_block_stmt_1873__entry__
      -- CP-element group 0: 	 branch_block_stmt_1873/do_while_stmt_1874__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1873/$exit
      -- CP-element group 1: 	 branch_block_stmt_1873/branch_block_stmt_1873__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1873/do_while_stmt_1874__exit__
      -- 
    timerDaemon_CP_3718_elements(1) <= timerDaemon_CP_3718_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1873/do_while_stmt_1874/$entry
      -- CP-element group 2: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874__entry__
      -- 
    timerDaemon_CP_3718_elements(2) <= timerDaemon_CP_3718_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874__exit__
      -- 
    -- Element group timerDaemon_CP_3718_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_back
      -- 
    -- Element group timerDaemon_CP_3718_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1873/do_while_stmt_1874/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_taken/$entry
      -- 
    timerDaemon_CP_3718_elements(5) <= timerDaemon_CP_3718_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_body_done
      -- 
    timerDaemon_CP_3718_elements(6) <= timerDaemon_CP_3718_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3718_elements(7) <= timerDaemon_CP_3718_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3718_elements(8) <= timerDaemon_CP_3718_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_3718_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/condition_evaluated
      -- 
    condition_evaluated_3742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(10), ack => do_while_stmt_1874_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(35) & timerDaemon_CP_3718_elements(15);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(12) & timerDaemon_CP_3718_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(9) & timerDaemon_CP_3718_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(9) & timerDaemon_CP_3718_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_3718_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_3718_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_loopback_trigger
      -- 
    timerDaemon_CP_3718_elements(16) <= timerDaemon_CP_3718_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_loopback_sample_req_ps
      -- 
    phi_stmt_1876_loopback_sample_req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1876_loopback_sample_req_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(17), ack => phi_stmt_1876_req_1); -- 
    -- Element group timerDaemon_CP_3718_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_entry_trigger
      -- 
    timerDaemon_CP_3718_elements(18) <= timerDaemon_CP_3718_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_entry_sample_req_ps
      -- 
    phi_stmt_1876_entry_sample_req_3760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1876_entry_sample_req_3760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(19), ack => phi_stmt_1876_req_0); -- 
    -- Element group timerDaemon_CP_3718_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/phi_stmt_1876_phi_mux_ack_ps
      -- 
    phi_stmt_1876_phi_mux_ack_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1876_ack_0, ack => timerDaemon_CP_3718_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_sample_completed_
      -- 
    -- Element group timerDaemon_CP_3718_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_update_start_
      -- 
    -- Element group timerDaemon_CP_3718_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_update_completed__ps
      -- 
    timerDaemon_CP_3718_elements(23) <= timerDaemon_CP_3718_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/type_cast_1879_update_completed_
      -- 
    -- Element group timerDaemon_CP_3718_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_3718_elements(22), ack => timerDaemon_CP_3718_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_3718_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_update_start__ps
      -- 
    -- Element group timerDaemon_CP_3718_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Sample/rr
      -- 
    rr_3784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(27), ack => ADD_u64_u64_1882_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(25) & timerDaemon_CP_3718_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Update/cr
      -- 
    cr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(28), ack => ADD_u64_u64_1882_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(26) & timerDaemon_CP_3718_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Sample/ra
      -- 
    ra_3785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1882_inst_ack_0, ack => timerDaemon_CP_3718_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/ADD_u64_u64_1882_Update/ca
      -- 
    ca_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1882_inst_ack_1, ack => timerDaemon_CP_3718_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/STORE_count_1884_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/STORE_count_1884_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/STORE_count_1884_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/STORE_count_1884_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/word_0/rr
      -- 
    rr_3812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(31), ack => STORE_count_1884_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(9) & timerDaemon_CP_3718_elements(15) & timerDaemon_CP_3718_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/word_0/cr
      -- 
    cr_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3718_elements(32), ack => STORE_count_1884_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_3718_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Sample/word_access_start/word_0/ra
      -- 
    ra_3813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1884_store_0_ack_0, ack => timerDaemon_CP_3718_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/STORE_count_1884_Update/word_access_complete/word_0/ca
      -- 
    ca_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1884_store_0_ack_1, ack => timerDaemon_CP_3718_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3718_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_3718_elements(9), ack => timerDaemon_CP_3718_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1873/do_while_stmt_1874/do_while_stmt_1874_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3718_elements(34) & timerDaemon_CP_3718_elements(14);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3718_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_exit/ack
      -- 
    ack_3829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1874_branch_ack_0, ack => timerDaemon_CP_3718_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_1873/do_while_stmt_1874/loop_taken/ack
      -- 
    ack_3833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1874_branch_ack_1, ack => timerDaemon_CP_3718_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1873/do_while_stmt_1874/$exit
      -- 
    timerDaemon_CP_3718_elements(39) <= timerDaemon_CP_3718_elements(3);
    timerDaemon_do_while_stmt_1874_terminator_3834: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1874_terminator_3834", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_3718_elements(6),loop_continue => timerDaemon_CP_3718_elements(38),loop_terminate => timerDaemon_CP_3718_elements(37),loop_back => timerDaemon_CP_3718_elements(4),loop_exit => timerDaemon_CP_3718_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1876_phi_seq_3791_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3718_elements(18);
      timerDaemon_CP_3718_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3718_elements(21);
      timerDaemon_CP_3718_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3718_elements(23);
      timerDaemon_CP_3718_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3718_elements(16);
      timerDaemon_CP_3718_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3718_elements(29);
      timerDaemon_CP_3718_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3718_elements(30);
      timerDaemon_CP_3718_elements(17) <= phi_mux_reqs(1);
      phi_stmt_1876_phi_seq_3791 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1876_phi_seq_3791") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3718_elements(11), 
          phi_sample_ack => timerDaemon_CP_3718_elements(14), 
          phi_update_req => timerDaemon_CP_3718_elements(13), 
          phi_update_ack => timerDaemon_CP_3718_elements(15), 
          phi_mux_ack => timerDaemon_CP_3718_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3743_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3718_elements(7);
        preds(1)  <= timerDaemon_CP_3718_elements(8);
        entry_tmerge_3743 : transition_merge -- 
          generic map(name => " entry_tmerge_3743")
          port map (preds => preds, symbol_out => timerDaemon_CP_3718_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_1882_wire : std_logic_vector(63 downto 0);
    signal STORE_count_1884_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_1884_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_1881_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1888_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_1876 : std_logic_vector(63 downto 0);
    signal type_cast_1879_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_1884_word_address_0 <= "0";
    konst_1881_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1888_wire_constant <= "1";
    type_cast_1879_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1876: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1879_wire_constant & ADD_u64_u64_1882_wire;
      req <= phi_stmt_1876_req_0 & phi_stmt_1876_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1876",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1876_ack_0,
          idata => idata,
          odata => ncount_1876,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1876
    -- equivalence STORE_count_1884_gather_scatter
    process(ncount_1876) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_1876;
      ov(63 downto 0) := iv;
      STORE_count_1884_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_1874_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1888_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1874_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1874_branch_req_0,
          ack0 => do_while_stmt_1874_branch_ack_0,
          ack1 => do_while_stmt_1874_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_1882_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_1876;
      ADD_u64_u64_1882_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1882_inst_req_0;
      ADD_u64_u64_1882_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1882_inst_req_1;
      ADD_u64_u64_1882_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_1884_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_1884_store_0_req_0;
      STORE_count_1884_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_1884_store_0_req_1;
      STORE_count_1884_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_1884_word_address_0;
      data_in <= STORE_count_1884_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module fill_T
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_T
  signal fill_T_addr :  std_logic_vector(63 downto 0);
  signal fill_T_in_args    : std_logic_vector(63 downto 0);
  signal fill_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_T_tag_out   : std_logic_vector(1 downto 0);
  signal fill_T_start_req : std_logic;
  signal fill_T_start_ack : std_logic;
  signal fill_T_fin_req   : std_logic;
  signal fill_T_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_T
  signal fill_T_call_reqs: std_logic_vector(0 downto 0);
  signal fill_T_call_acks: std_logic_vector(0 downto 0);
  signal fill_T_return_reqs: std_logic_vector(0 downto 0);
  signal fill_T_return_acks: std_logic_vector(0 downto 0);
  signal fill_T_call_data: std_logic_vector(63 downto 0);
  signal fill_T_call_tag: std_logic_vector(0 downto 0);
  signal fill_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool3D
  component maxPool3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(159 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool3D
  signal maxPool3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool3D_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool3D_start_req : std_logic;
  signal maxPool3D_start_ack : std_logic;
  signal maxPool3D_fin_req   : std_logic;
  signal maxPool3D_fin_ack : std_logic;
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(159 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(159 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_T
  fill_T_addr <= fill_T_in_args(63 downto 0);
  -- call arbiter for module fill_T
  fill_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_T_call_reqs,
      call_acks => fill_T_call_acks,
      return_reqs => fill_T_return_reqs,
      return_acks => fill_T_return_acks,
      call_data  => fill_T_call_data,
      call_tag  => fill_T_call_tag,
      return_tag  => fill_T_return_tag,
      call_mtag => fill_T_tag_in,
      return_mtag => fill_T_tag_out,
      call_mreq => fill_T_start_req,
      call_mack => fill_T_start_ack,
      return_mreq => fill_T_fin_req,
      return_mack => fill_T_fin_ack,
      call_mdata => fill_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_T_instance:fill_T-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_T_addr,
      start_req => fill_T_start_req,
      start_ack => fill_T_start_ack,
      fin_req => fill_T_fin_req,
      fin_ack => fill_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(255 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(1 downto 1),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(1 downto 1),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 8),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => fill_T_tag_in,
      tag_out => fill_T_tag_out-- 
    ); -- 
  -- module maxPool3D
  maxPool3D_instance:maxPool3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => maxPool3D_start_req,
      start_ack => maxPool3D_start_ack,
      fin_req => maxPool3D_fin_req,
      fin_ack => maxPool3D_fin_ack,
      clk => clk,
      reset => reset,
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      fill_T_call_reqs => fill_T_call_reqs(0 downto 0),
      fill_T_call_acks => fill_T_call_acks(0 downto 0),
      fill_T_call_data => fill_T_call_data(63 downto 0),
      fill_T_call_tag => fill_T_call_tag(0 downto 0),
      fill_T_return_reqs => fill_T_return_reqs(0 downto 0),
      fill_T_return_acks => fill_T_return_acks(0 downto 0),
      fill_T_return_tag => fill_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(159 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => maxPool3D_tag_in,
      tag_out => maxPool3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  maxPool3D_tag_in <= (others => '0');
  maxPool3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => maxPool3D_start_req, start_ack => maxPool3D_start_ack,  fin_req => maxPool3D_fin_req,  fin_ack => maxPool3D_fin_ack);
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(159 downto 128);
  maxPool4_addr1 <= maxPool4_in_args(127 downto 96);
  maxPool4_addr2 <= maxPool4_in_args(95 downto 64);
  maxPool4_addr3 <= maxPool4_in_args(63 downto 32);
  maxPool4_addr4 <= maxPool4_in_args(31 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 160,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 256,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 256
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
