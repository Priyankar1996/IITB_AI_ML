-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3648_start: Boolean;
  signal convTranspose_CP_3648_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1227_call_req_0 : boolean;
  signal call_stmt_1227_call_ack_0 : boolean;
  signal call_stmt_1227_call_req_1 : boolean;
  signal call_stmt_1227_call_ack_1 : boolean;
  signal WPIPE_Block0_start_1229_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1229_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1229_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1229_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1232_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1232_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1232_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1232_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1235_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1235_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1235_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1235_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1238_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1238_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1238_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1238_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1243_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1243_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1243_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1243_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1246_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1246_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1246_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1246_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1249_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1249_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1249_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1249_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1252_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1252_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1252_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1252_inst_ack_1 : boolean;
  signal call_stmt_1255_call_req_0 : boolean;
  signal call_stmt_1255_call_ack_0 : boolean;
  signal call_stmt_1255_call_req_1 : boolean;
  signal call_stmt_1255_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3648_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3648_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3648_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3648_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3648: Block -- control-path 
    signal convTranspose_CP_3648_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3648_elements(0) <= convTranspose_CP_3648_start;
    convTranspose_CP_3648_symbol <= convTranspose_CP_3648_elements(22);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1225/$entry
      -- CP-element group 0: 	 branch_block_stmt_1225/branch_block_stmt_1225__entry__
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227__entry__
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/$entry
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Update/ccr
      -- 
    crr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(0), ack => call_stmt_1227_call_req_0); -- 
    ccr_3681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(0), ack => call_stmt_1227_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Sample/cra
      -- 
    cra_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1227_call_ack_0, ack => convTranspose_CP_3648_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (19) 
      -- CP-element group 2: 	 branch_block_stmt_1225/call_stmt_1227__exit__
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240__entry__
      -- CP-element group 2: 	 branch_block_stmt_1225/call_stmt_1227/$exit
      -- CP-element group 2: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1225/call_stmt_1227/call_stmt_1227_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/$entry
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Sample/req
      -- 
    cca_3682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1227_call_ack_1, ack => convTranspose_CP_3648_elements(2)); -- 
    req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(2), ack => WPIPE_Block0_start_1229_inst_req_0); -- 
    req_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(2), ack => WPIPE_Block1_start_1232_inst_req_0); -- 
    req_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(2), ack => WPIPE_Block2_start_1235_inst_req_0); -- 
    req_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(2), ack => WPIPE_Block3_start_1238_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Update/req
      -- 
    ack_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1229_inst_ack_0, ack => convTranspose_CP_3648_elements(3)); -- 
    req_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(3), ack => WPIPE_Block0_start_1229_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block0_start_1229_Update/ack
      -- 
    ack_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1229_inst_ack_1, ack => convTranspose_CP_3648_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Update/req
      -- 
    ack_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1232_inst_ack_0, ack => convTranspose_CP_3648_elements(5)); -- 
    req_3712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(5), ack => WPIPE_Block1_start_1232_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	11 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block1_start_1232_Update/ack
      -- 
    ack_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1232_inst_ack_1, ack => convTranspose_CP_3648_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Update/req
      -- 
    ack_3722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1235_inst_ack_0, ack => convTranspose_CP_3648_elements(7)); -- 
    req_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(7), ack => WPIPE_Block2_start_1235_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block2_start_1235_Update/ack
      -- 
    ack_3727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1235_inst_ack_1, ack => convTranspose_CP_3648_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Update/req
      -- 
    ack_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1238_inst_ack_0, ack => convTranspose_CP_3648_elements(9)); -- 
    req_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(9), ack => WPIPE_Block3_start_1238_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/WPIPE_Block3_start_1238_Update/ack
      -- 
    ack_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1238_inst_ack_1, ack => convTranspose_CP_3648_elements(10)); -- 
    -- CP-element group 11:  join  fork  transition  place  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	6 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240__exit__
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253__entry__
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1231_to_assign_stmt_1240/$exit
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/$entry
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Sample/rr
      -- 
    rr_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(11), ack => RPIPE_Block0_done_1243_inst_req_0); -- 
    rr_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(11), ack => RPIPE_Block1_done_1246_inst_req_0); -- 
    rr_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(11), ack => RPIPE_Block2_done_1249_inst_req_0); -- 
    rr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(11), ack => RPIPE_Block3_done_1252_inst_req_0); -- 
    convTranspose_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_3648_elements(8) & convTranspose_CP_3648_elements(4) & convTranspose_CP_3648_elements(10) & convTranspose_CP_3648_elements(6);
      gj_convTranspose_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3648_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Update/cr
      -- 
    ra_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1243_inst_ack_0, ack => convTranspose_CP_3648_elements(12)); -- 
    cr_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(12), ack => RPIPE_Block0_done_1243_inst_req_1); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block0_done_1243_Update/ca
      -- 
    ca_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1243_inst_ack_1, ack => convTranspose_CP_3648_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Update/cr
      -- 
    ra_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1246_inst_ack_0, ack => convTranspose_CP_3648_elements(14)); -- 
    cr_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(14), ack => RPIPE_Block1_done_1246_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block1_done_1246_Update/ca
      -- 
    ca_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1246_inst_ack_1, ack => convTranspose_CP_3648_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Update/cr
      -- 
    ra_3781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1249_inst_ack_0, ack => convTranspose_CP_3648_elements(16)); -- 
    cr_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(16), ack => RPIPE_Block2_done_1249_inst_req_1); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block2_done_1249_Update/ca
      -- 
    ca_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1249_inst_ack_1, ack => convTranspose_CP_3648_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Update/cr
      -- 
    ra_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1252_inst_ack_0, ack => convTranspose_CP_3648_elements(18)); -- 
    cr_3799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(18), ack => RPIPE_Block3_done_1252_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/RPIPE_Block3_done_1252_Update/ca
      -- 
    ca_3800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1252_inst_ack_1, ack => convTranspose_CP_3648_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  place  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	13 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (10) 
      -- CP-element group 20: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253__exit__
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255__entry__
      -- CP-element group 20: 	 branch_block_stmt_1225/assign_stmt_1244_to_assign_stmt_1253/$exit
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/$entry
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Sample/crr
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Update/ccr
      -- 
    crr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(20), ack => call_stmt_1255_call_req_0); -- 
    ccr_3816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3648_elements(20), ack => call_stmt_1255_call_req_1); -- 
    convTranspose_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_3648_elements(13) & convTranspose_CP_3648_elements(17) & convTranspose_CP_3648_elements(15) & convTranspose_CP_3648_elements(19);
      gj_convTranspose_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3648_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Sample/cra
      -- 
    cra_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1255_call_ack_0, ack => convTranspose_CP_3648_elements(21)); -- 
    -- CP-element group 22:  transition  place  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (16) 
      -- CP-element group 22: 	 $exit
      -- CP-element group 22: 	 branch_block_stmt_1225/$exit
      -- CP-element group 22: 	 branch_block_stmt_1225/branch_block_stmt_1225__exit__
      -- CP-element group 22: 	 branch_block_stmt_1225/call_stmt_1255__exit__
      -- CP-element group 22: 	 branch_block_stmt_1225/return__
      -- CP-element group 22: 	 branch_block_stmt_1225/merge_stmt_1257__exit__
      -- CP-element group 22: 	 branch_block_stmt_1225/call_stmt_1255/$exit
      -- CP-element group 22: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1225/call_stmt_1255/call_stmt_1255_Update/cca
      -- CP-element group 22: 	 branch_block_stmt_1225/return___PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_1225/return___PhiReq/$exit
      -- CP-element group 22: 	 branch_block_stmt_1225/merge_stmt_1257_PhiReqMerge
      -- CP-element group 22: 	 branch_block_stmt_1225/merge_stmt_1257_PhiAck/$entry
      -- CP-element group 22: 	 branch_block_stmt_1225/merge_stmt_1257_PhiAck/$exit
      -- CP-element group 22: 	 branch_block_stmt_1225/merge_stmt_1257_PhiAck/dummy
      -- 
    cca_3817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1255_call_ack_1, ack => convTranspose_CP_3648_elements(22)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call11_1253 : std_logic_vector(15 downto 0);
    signal call5_1244 : std_logic_vector(15 downto 0);
    signal call7_1247 : std_logic_vector(15 downto 0);
    signal call9_1250 : std_logic_vector(15 downto 0);
    signal call_1227 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- shared inport operator group (0) : RPIPE_Block0_done_1243_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1243_inst_req_0;
      RPIPE_Block0_done_1243_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1243_inst_req_1;
      RPIPE_Block0_done_1243_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call5_1244 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1246_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1246_inst_req_0;
      RPIPE_Block1_done_1246_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1246_inst_req_1;
      RPIPE_Block1_done_1246_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call7_1247 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1249_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1249_inst_req_0;
      RPIPE_Block2_done_1249_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1249_inst_req_1;
      RPIPE_Block2_done_1249_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call9_1250 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1252_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1252_inst_req_0;
      RPIPE_Block3_done_1252_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1252_inst_req_1;
      RPIPE_Block3_done_1252_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call11_1253 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1229_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1229_inst_req_0;
      WPIPE_Block0_start_1229_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1229_inst_req_1;
      WPIPE_Block0_start_1229_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1227;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1232_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1232_inst_req_0;
      WPIPE_Block1_start_1232_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1232_inst_req_1;
      WPIPE_Block1_start_1232_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1227;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1235_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1235_inst_req_0;
      WPIPE_Block2_start_1235_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1235_inst_req_1;
      WPIPE_Block2_start_1235_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1227;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1238_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1238_inst_req_0;
      WPIPE_Block3_start_1238_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1238_inst_req_1;
      WPIPE_Block3_start_1238_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1227;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1227_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1227_call_req_0;
      call_stmt_1227_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1227_call_req_1;
      call_stmt_1227_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1227 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1255_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1255_call_req_0;
      call_stmt_1255_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1255_call_req_1;
      call_stmt_1255_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3826_start: Boolean;
  signal convTransposeA_CP_3826_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1298_load_0_req_0 : boolean;
  signal RPIPE_Block0_start_1263_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1263_inst_ack_0 : boolean;
  signal ptr_deref_1288_load_0_req_1 : boolean;
  signal RPIPE_Block0_start_1263_inst_req_1 : boolean;
  signal ptr_deref_1298_load_0_ack_0 : boolean;
  signal ptr_deref_1288_load_0_ack_1 : boolean;
  signal ptr_deref_1288_load_0_req_0 : boolean;
  signal RPIPE_Block0_start_1263_inst_ack_1 : boolean;
  signal ptr_deref_1288_load_0_ack_0 : boolean;
  signal LOAD_padding_1313_load_0_req_1 : boolean;
  signal LOAD_padding_1313_load_0_ack_1 : boolean;
  signal ptr_deref_1276_load_0_ack_1 : boolean;
  signal ptr_deref_1276_load_0_req_1 : boolean;
  signal LOAD_padding_1313_load_0_req_0 : boolean;
  signal LOAD_padding_1313_load_0_ack_0 : boolean;
  signal ptr_deref_1310_load_0_req_0 : boolean;
  signal ptr_deref_1310_load_0_ack_0 : boolean;
  signal ptr_deref_1310_load_0_req_1 : boolean;
  signal ptr_deref_1310_load_0_ack_1 : boolean;
  signal ptr_deref_1276_load_0_ack_0 : boolean;
  signal ptr_deref_1298_load_0_ack_1 : boolean;
  signal ptr_deref_1276_load_0_req_0 : boolean;
  signal ptr_deref_1298_load_0_req_1 : boolean;
  signal ptr_deref_1323_load_0_req_0 : boolean;
  signal ptr_deref_1323_load_0_ack_0 : boolean;
  signal ptr_deref_1323_load_0_req_1 : boolean;
  signal ptr_deref_1323_load_0_ack_1 : boolean;
  signal ptr_deref_1335_load_0_req_0 : boolean;
  signal ptr_deref_1335_load_0_ack_0 : boolean;
  signal ptr_deref_1335_load_0_req_1 : boolean;
  signal ptr_deref_1335_load_0_ack_1 : boolean;
  signal ptr_deref_1347_load_0_req_0 : boolean;
  signal ptr_deref_1347_load_0_ack_0 : boolean;
  signal ptr_deref_1347_load_0_req_1 : boolean;
  signal ptr_deref_1347_load_0_ack_1 : boolean;
  signal ptr_deref_1359_load_0_req_0 : boolean;
  signal ptr_deref_1359_load_0_ack_0 : boolean;
  signal ptr_deref_1359_load_0_req_1 : boolean;
  signal ptr_deref_1359_load_0_ack_1 : boolean;
  signal type_cast_1363_inst_req_0 : boolean;
  signal type_cast_1363_inst_ack_0 : boolean;
  signal type_cast_1363_inst_req_1 : boolean;
  signal type_cast_1363_inst_ack_1 : boolean;
  signal type_cast_1367_inst_req_0 : boolean;
  signal type_cast_1367_inst_ack_0 : boolean;
  signal type_cast_1367_inst_req_1 : boolean;
  signal type_cast_1367_inst_ack_1 : boolean;
  signal ptr_deref_1385_load_0_req_0 : boolean;
  signal ptr_deref_1385_load_0_ack_0 : boolean;
  signal ptr_deref_1385_load_0_req_1 : boolean;
  signal ptr_deref_1385_load_0_ack_1 : boolean;
  signal type_cast_1389_inst_req_0 : boolean;
  signal type_cast_1389_inst_ack_0 : boolean;
  signal type_cast_1389_inst_req_1 : boolean;
  signal type_cast_1389_inst_ack_1 : boolean;
  signal type_cast_1514_inst_req_0 : boolean;
  signal type_cast_1514_inst_ack_0 : boolean;
  signal type_cast_1514_inst_req_1 : boolean;
  signal type_cast_1514_inst_ack_1 : boolean;
  signal array_obj_ref_1526_index_offset_req_0 : boolean;
  signal array_obj_ref_1526_index_offset_ack_0 : boolean;
  signal array_obj_ref_1526_index_offset_req_1 : boolean;
  signal array_obj_ref_1526_index_offset_ack_1 : boolean;
  signal addr_of_1527_final_reg_req_0 : boolean;
  signal addr_of_1527_final_reg_ack_0 : boolean;
  signal addr_of_1527_final_reg_req_1 : boolean;
  signal addr_of_1527_final_reg_ack_1 : boolean;
  signal ptr_deref_1531_load_0_req_0 : boolean;
  signal ptr_deref_1531_load_0_ack_0 : boolean;
  signal ptr_deref_1531_load_0_req_1 : boolean;
  signal ptr_deref_1531_load_0_ack_1 : boolean;
  signal type_cast_1535_inst_req_0 : boolean;
  signal type_cast_1535_inst_ack_0 : boolean;
  signal type_cast_1535_inst_req_1 : boolean;
  signal type_cast_1535_inst_ack_1 : boolean;
  signal array_obj_ref_1547_index_offset_req_0 : boolean;
  signal array_obj_ref_1547_index_offset_ack_0 : boolean;
  signal array_obj_ref_1547_index_offset_req_1 : boolean;
  signal array_obj_ref_1547_index_offset_ack_1 : boolean;
  signal addr_of_1548_final_reg_req_0 : boolean;
  signal addr_of_1548_final_reg_ack_0 : boolean;
  signal addr_of_1548_final_reg_req_1 : boolean;
  signal addr_of_1548_final_reg_ack_1 : boolean;
  signal ptr_deref_1551_store_0_req_0 : boolean;
  signal ptr_deref_1551_store_0_ack_0 : boolean;
  signal ptr_deref_1551_store_0_req_1 : boolean;
  signal ptr_deref_1551_store_0_ack_1 : boolean;
  signal type_cast_1556_inst_req_0 : boolean;
  signal type_cast_1556_inst_ack_0 : boolean;
  signal type_cast_1556_inst_req_1 : boolean;
  signal type_cast_1556_inst_ack_1 : boolean;
  signal if_stmt_1569_branch_req_0 : boolean;
  signal if_stmt_1569_branch_ack_1 : boolean;
  signal if_stmt_1569_branch_ack_0 : boolean;
  signal type_cast_1592_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_0 : boolean;
  signal type_cast_1592_inst_req_1 : boolean;
  signal type_cast_1592_inst_ack_1 : boolean;
  signal type_cast_1601_inst_req_0 : boolean;
  signal type_cast_1601_inst_ack_0 : boolean;
  signal type_cast_1601_inst_req_1 : boolean;
  signal type_cast_1601_inst_ack_1 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_1 : boolean;
  signal type_cast_1617_inst_ack_1 : boolean;
  signal if_stmt_1624_branch_req_0 : boolean;
  signal if_stmt_1624_branch_ack_1 : boolean;
  signal if_stmt_1624_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1632_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1632_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1632_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1632_inst_ack_1 : boolean;
  signal phi_stmt_1421_req_0 : boolean;
  signal phi_stmt_1428_req_0 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal type_cast_1427_inst_req_1 : boolean;
  signal type_cast_1427_inst_ack_1 : boolean;
  signal phi_stmt_1421_req_1 : boolean;
  signal type_cast_1434_inst_req_0 : boolean;
  signal type_cast_1434_inst_ack_0 : boolean;
  signal type_cast_1434_inst_req_1 : boolean;
  signal type_cast_1434_inst_ack_1 : boolean;
  signal phi_stmt_1428_req_1 : boolean;
  signal phi_stmt_1421_ack_0 : boolean;
  signal phi_stmt_1428_ack_0 : boolean;
  signal type_cast_1494_inst_req_0 : boolean;
  signal type_cast_1494_inst_ack_0 : boolean;
  signal type_cast_1494_inst_req_1 : boolean;
  signal type_cast_1494_inst_ack_1 : boolean;
  signal phi_stmt_1488_req_1 : boolean;
  signal phi_stmt_1488_req_0 : boolean;
  signal phi_stmt_1488_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3826_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3826_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3826_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3826_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3826: Block -- control-path 
    signal convTransposeA_CP_3826_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3826_elements(0) <= convTransposeA_CP_3826_start;
    convTransposeA_CP_3826_symbol <= convTransposeA_CP_3826_elements(61);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1261/assign_stmt_1264/$entry
      -- CP-element group 0: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1261/assign_stmt_1264__entry__
      -- CP-element group 0: 	 branch_block_stmt_1261/branch_block_stmt_1261__entry__
      -- CP-element group 0: 	 branch_block_stmt_1261/$entry
      -- CP-element group 0: 	 $entry
      -- 
    rr_3874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(0), ack => RPIPE_Block0_start_1263_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Update/$entry
      -- 
    ra_3875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1263_inst_ack_0, ack => convTransposeA_CP_3826_elements(1)); -- 
    cr_3879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(1), ack => RPIPE_Block0_start_1263_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1264/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1264__exit__
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418__entry__
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1264/RPIPE_Block0_start_1263_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Update/cr
      -- 
    ca_3880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1263_inst_ack_1, ack => convTransposeA_CP_3826_elements(2)); -- 
    rr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1298_load_0_req_0); -- 
    cr_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1288_load_0_req_1); -- 
    rr_3966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1288_load_0_req_0); -- 
    cr_4110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => LOAD_padding_1313_load_0_req_1); -- 
    cr_3927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1276_load_0_req_1); -- 
    rr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => LOAD_padding_1313_load_0_req_0); -- 
    rr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1310_load_0_req_0); -- 
    cr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1310_load_0_req_1); -- 
    rr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1276_load_0_req_0); -- 
    cr_4027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1298_load_0_req_1); -- 
    rr_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1323_load_0_req_0); -- 
    cr_4160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1323_load_0_req_1); -- 
    rr_4199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1335_load_0_req_0); -- 
    cr_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1335_load_0_req_1); -- 
    rr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1347_load_0_req_0); -- 
    cr_4260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1347_load_0_req_1); -- 
    rr_4299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1359_load_0_req_0); -- 
    cr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1359_load_0_req_1); -- 
    cr_4329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => type_cast_1363_inst_req_1); -- 
    cr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => type_cast_1367_inst_req_1); -- 
    rr_4377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1385_load_0_req_0); -- 
    cr_4388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => ptr_deref_1385_load_0_req_1); -- 
    cr_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(2), ack => type_cast_1389_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Sample/word_access_start/word_0/$exit
      -- 
    ra_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1276_load_0_ack_0, ack => convTransposeA_CP_3826_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	21 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/ptr_deref_1276_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/ptr_deref_1276_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/ptr_deref_1276_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/ptr_deref_1276_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1276_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Sample/rr
      -- 
    ca_3928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1276_load_0_ack_1, ack => convTransposeA_CP_3826_elements(4)); -- 
    rr_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(4), ack => type_cast_1363_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Sample/word_access_start/word_0/ra
      -- 
    ra_3967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1288_load_0_ack_0, ack => convTransposeA_CP_3826_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/ptr_deref_1288_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/ptr_deref_1288_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/ptr_deref_1288_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1288_Update/ptr_deref_1288_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Sample/rr
      -- 
    ca_3978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1288_load_0_ack_1, ack => convTransposeA_CP_3826_elements(6)); -- 
    rr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(6), ack => type_cast_1367_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Sample/$exit
      -- 
    ra_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1298_load_0_ack_0, ack => convTransposeA_CP_3826_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	29 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/ptr_deref_1298_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/ptr_deref_1298_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/ptr_deref_1298_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/ptr_deref_1298_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1298_Update/word_access_complete/word_0/ca
      -- 
    ca_4028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1298_load_0_ack_1, ack => convTransposeA_CP_3826_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Sample/word_access_start/word_0/$exit
      -- 
    ra_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1310_load_0_ack_0, ack => convTransposeA_CP_3826_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/ptr_deref_1310_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/ptr_deref_1310_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/ptr_deref_1310_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1310_Update/ptr_deref_1310_Merge/merge_ack
      -- 
    ca_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1310_load_0_ack_1, ack => convTransposeA_CP_3826_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Sample/word_access_start/word_0/ra
      -- 
    ra_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1313_load_0_ack_0, ack => convTransposeA_CP_3826_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/LOAD_padding_1313_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/LOAD_padding_1313_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/LOAD_padding_1313_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_Update/LOAD_padding_1313_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/LOAD_padding_1313_update_completed_
      -- 
    ca_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1313_load_0_ack_1, ack => convTransposeA_CP_3826_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Sample/word_access_start/word_0/ra
      -- 
    ra_4150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1323_load_0_ack_0, ack => convTransposeA_CP_3826_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/ptr_deref_1323_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/ptr_deref_1323_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/ptr_deref_1323_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1323_Update/ptr_deref_1323_Merge/merge_ack
      -- 
    ca_4161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1323_load_0_ack_1, ack => convTransposeA_CP_3826_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Sample/word_access_start/word_0/ra
      -- 
    ra_4200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1335_load_0_ack_0, ack => convTransposeA_CP_3826_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/ptr_deref_1335_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/ptr_deref_1335_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/ptr_deref_1335_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1335_Update/ptr_deref_1335_Merge/merge_ack
      -- 
    ca_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1335_load_0_ack_1, ack => convTransposeA_CP_3826_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Sample/word_access_start/word_0/ra
      -- 
    ra_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1347_load_0_ack_0, ack => convTransposeA_CP_3826_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/ptr_deref_1347_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/ptr_deref_1347_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/ptr_deref_1347_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1347_Update/ptr_deref_1347_Merge/merge_ack
      -- 
    ca_4261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1347_load_0_ack_1, ack => convTransposeA_CP_3826_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Sample/word_access_start/word_0/ra
      -- 
    ra_4300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1359_load_0_ack_0, ack => convTransposeA_CP_3826_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/ptr_deref_1359_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/ptr_deref_1359_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/ptr_deref_1359_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1359_Update/ptr_deref_1359_Merge/merge_ack
      -- 
    ca_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1359_load_0_ack_1, ack => convTransposeA_CP_3826_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	4 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Sample/ra
      -- 
    ra_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_0, ack => convTransposeA_CP_3826_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1363_Update/ca
      -- 
    ca_4330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_1, ack => convTransposeA_CP_3826_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Sample/ra
      -- 
    ra_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1367_inst_ack_0, ack => convTransposeA_CP_3826_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1367_Update/ca
      -- 
    ca_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1367_inst_ack_1, ack => convTransposeA_CP_3826_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Sample/word_access_start/word_0/ra
      -- 
    ra_4378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1385_load_0_ack_0, ack => convTransposeA_CP_3826_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (12) 
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/ptr_deref_1385_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/ptr_deref_1385_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/ptr_deref_1385_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/ptr_deref_1385_Update/ptr_deref_1385_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Sample/rr
      -- 
    ca_4389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1385_load_0_ack_1, ack => convTransposeA_CP_3826_elements(26)); -- 
    rr_4402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(26), ack => type_cast_1389_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Sample/ra
      -- 
    ra_4403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_0, ack => convTransposeA_CP_3826_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/type_cast_1389_Update/ca
      -- 
    ca_4408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_1, ack => convTransposeA_CP_3826_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	8 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	14 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	62 
    -- CP-element group 29: 	63 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418__exit__
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1261/assign_stmt_1273_to_assign_stmt_1418/$exit
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/$entry
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/$entry
      -- CP-element group 29: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(8) & convTransposeA_CP_3826_elements(10) & convTransposeA_CP_3826_elements(12) & convTransposeA_CP_3826_elements(14) & convTransposeA_CP_3826_elements(16) & convTransposeA_CP_3826_elements(18) & convTransposeA_CP_3826_elements(20) & convTransposeA_CP_3826_elements(22) & convTransposeA_CP_3826_elements(24) & convTransposeA_CP_3826_elements(28);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	81 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Sample/ra
      -- 
    ra_4423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1514_inst_ack_0, ack => convTransposeA_CP_3826_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	81 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (16) 
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_resized_1
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_scaled_1
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_computed_1
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_resize_1/$entry
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_resize_1/$exit
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_resize_1/index_resize_req
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_resize_1/index_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_scale_1/$entry
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_scale_1/$exit
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_scale_1/scale_rename_req
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_index_scale_1/scale_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Sample/req
      -- 
    ca_4428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1514_inst_ack_1, ack => convTransposeA_CP_3826_elements(31)); -- 
    req_4453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(31), ack => array_obj_ref_1526_index_offset_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	49 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Sample/ack
      -- 
    ack_4454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1526_index_offset_ack_0, ack => convTransposeA_CP_3826_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	81 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (11) 
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_offset_calculated
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_request/$entry
      -- CP-element group 33: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_request/req
      -- 
    ack_4459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1526_index_offset_ack_1, ack => convTransposeA_CP_3826_elements(33)); -- 
    req_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(33), ack => addr_of_1527_final_reg_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_request/$exit
      -- CP-element group 34: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_request/ack
      -- 
    ack_4469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1527_final_reg_ack_0, ack => convTransposeA_CP_3826_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	81 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (24) 
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_complete/ack
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_word_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_address_resized
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_addr_resize/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_addr_resize/$exit
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_word_addrgen/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_word_addrgen/$exit
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_word_addrgen/root_register_req
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_word_addrgen/root_register_ack
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/word_0/rr
      -- 
    ack_4474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1527_final_reg_ack_1, ack => convTransposeA_CP_3826_elements(35)); -- 
    rr_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(35), ack => ptr_deref_1531_load_0_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Sample/word_access_start/word_0/ra
      -- 
    ra_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1531_load_0_ack_0, ack => convTransposeA_CP_3826_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	81 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	44 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/ptr_deref_1531_Merge/$entry
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/ptr_deref_1531_Merge/$exit
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/ptr_deref_1531_Merge/merge_req
      -- CP-element group 37: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/ptr_deref_1531_Merge/merge_ack
      -- 
    ca_4519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1531_load_0_ack_1, ack => convTransposeA_CP_3826_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	81 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Sample/ra
      -- 
    ra_4533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_0, ack => convTransposeA_CP_3826_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	81 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (16) 
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_resized_1
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_scaled_1
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_computed_1
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_resize_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_resize_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_resize_1/index_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_resize_1/index_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_scale_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_scale_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_scale_1/scale_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_index_scale_1/scale_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Sample/req
      -- 
    ca_4538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1535_inst_ack_1, ack => convTransposeA_CP_3826_elements(39)); -- 
    req_4563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(39), ack => array_obj_ref_1547_index_offset_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Sample/ack
      -- 
    ack_4564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1547_index_offset_ack_0, ack => convTransposeA_CP_3826_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	81 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_request/req
      -- 
    ack_4569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1547_index_offset_ack_1, ack => convTransposeA_CP_3826_elements(41)); -- 
    req_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(41), ack => addr_of_1548_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_request/ack
      -- 
    ack_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1548_final_reg_ack_0, ack => convTransposeA_CP_3826_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	81 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_word_addrgen/root_register_ack
      -- 
    ack_4584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1548_final_reg_ack_1, ack => convTransposeA_CP_3826_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	37 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/ptr_deref_1551_Split/$entry
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/ptr_deref_1551_Split/$exit
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_req
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/ptr_deref_1551_Split/split_ack
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/word_0/rr
      -- 
    rr_4622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(44), ack => ptr_deref_1551_store_0_req_0); -- 
    convTransposeA_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(37) & convTransposeA_CP_3826_elements(43);
      gj_convTransposeA_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Sample/word_access_start/word_0/ra
      -- 
    ra_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_0, ack => convTransposeA_CP_3826_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	81 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/word_0/ca
      -- 
    ca_4634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1551_store_0_ack_1, ack => convTransposeA_CP_3826_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	81 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Sample/ra
      -- 
    ra_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1556_inst_ack_0, ack => convTransposeA_CP_3826_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	81 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Update/ca
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1556_inst_ack_1, ack => convTransposeA_CP_3826_elements(48)); -- 
    -- CP-element group 49:  branch  join  transition  place  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	32 
    -- CP-element group 49: 	40 
    -- CP-element group 49: 	46 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (10) 
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569__entry__
      -- CP-element group 49: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568__exit__
      -- CP-element group 49: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/$exit
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_dead_link/$entry
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_eval_test/$entry
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_eval_test/$exit
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_eval_test/branch_req
      -- CP-element group 49: 	 branch_block_stmt_1261/R_cmp_1570_place
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_if_link/$entry
      -- CP-element group 49: 	 branch_block_stmt_1261/if_stmt_1569_else_link/$entry
      -- 
    branch_req_4656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(49), ack => if_stmt_1569_branch_req_0); -- 
    convTransposeA_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(32) & convTransposeA_CP_3826_elements(40) & convTransposeA_CP_3826_elements(46) & convTransposeA_CP_3826_elements(48);
      gj_convTransposeA_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	76 
    -- CP-element group 50: 	77 
    -- CP-element group 50:  members (24) 
      -- CP-element group 50: 	 branch_block_stmt_1261/assign_stmt_1581__exit__
      -- CP-element group 50: 	 branch_block_stmt_1261/assign_stmt_1581__entry__
      -- CP-element group 50: 	 branch_block_stmt_1261/merge_stmt_1575__exit__
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody
      -- CP-element group 50: 	 branch_block_stmt_1261/if_stmt_1569_if_link/$exit
      -- CP-element group 50: 	 branch_block_stmt_1261/if_stmt_1569_if_link/if_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_1261/whilex_xbody_ifx_xthen
      -- CP-element group 50: 	 branch_block_stmt_1261/assign_stmt_1581/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/assign_stmt_1581/$exit
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1261/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 50: 	 branch_block_stmt_1261/merge_stmt_1575_PhiReqMerge
      -- CP-element group 50: 	 branch_block_stmt_1261/merge_stmt_1575_PhiAck/$entry
      -- CP-element group 50: 	 branch_block_stmt_1261/merge_stmt_1575_PhiAck/$exit
      -- CP-element group 50: 	 branch_block_stmt_1261/merge_stmt_1575_PhiAck/dummy
      -- 
    if_choice_transition_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1569_branch_ack_1, ack => convTransposeA_CP_3826_elements(50)); -- 
    rr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(50), ack => type_cast_1494_inst_req_0); -- 
    cr_4849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(50), ack => type_cast_1494_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	55 
    -- CP-element group 51: 	57 
    -- CP-element group 51:  members (24) 
      -- CP-element group 51: 	 branch_block_stmt_1261/merge_stmt_1583__exit__
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623__entry__
      -- CP-element group 51: 	 branch_block_stmt_1261/merge_stmt_1583_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_1261/merge_stmt_1583_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_1261/merge_stmt_1583_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1261/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/merge_stmt_1583_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_1261/if_stmt_1569_else_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1261/if_stmt_1569_else_link/else_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1261/whilex_xbody_ifx_xelse
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Update/cr
      -- 
    else_choice_transition_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1569_branch_ack_0, ack => convTransposeA_CP_3826_elements(51)); -- 
    rr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(51), ack => type_cast_1592_inst_req_0); -- 
    cr_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(51), ack => type_cast_1592_inst_req_1); -- 
    cr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(51), ack => type_cast_1601_inst_req_1); -- 
    cr_4714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(51), ack => type_cast_1617_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Sample/ra
      -- 
    ra_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_0, ack => convTransposeA_CP_3826_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1592_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Sample/rr
      -- 
    ca_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_1, ack => convTransposeA_CP_3826_elements(53)); -- 
    rr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(53), ack => type_cast_1601_inst_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Sample/ra
      -- 
    ra_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_0, ack => convTransposeA_CP_3826_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	51 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1601_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Sample/rr
      -- 
    ca_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1601_inst_ack_1, ack => convTransposeA_CP_3826_elements(55)); -- 
    rr_4709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(55), ack => type_cast_1617_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Sample/ra
      -- 
    ra_4710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_0, ack => convTransposeA_CP_3826_elements(56)); -- 
    -- CP-element group 57:  branch  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623__exit__
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624__entry__
      -- CP-element group 57: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/$exit
      -- CP-element group 57: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1261/assign_stmt_1589_to_assign_stmt_1623/type_cast_1617_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1261/R_cmp86_1625_place
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1261/if_stmt_1624_else_link/$entry
      -- 
    ca_4715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_1, ack => convTransposeA_CP_3826_elements(57)); -- 
    branch_req_4723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(57), ack => if_stmt_1624_branch_req_0); -- 
    -- CP-element group 58:  merge  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (15) 
      -- CP-element group 58: 	 branch_block_stmt_1261/merge_stmt_1630__exit__
      -- CP-element group 58: 	 branch_block_stmt_1261/assign_stmt_1634__entry__
      -- CP-element group 58: 	 branch_block_stmt_1261/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1261/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1261/merge_stmt_1630_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1261/merge_stmt_1630_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1261/merge_stmt_1630_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1261/merge_stmt_1630_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1261/if_stmt_1624_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1261/if_stmt_1624_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1261/ifx_xelse_whilex_xend
      -- CP-element group 58: 	 branch_block_stmt_1261/assign_stmt_1634/$entry
      -- CP-element group 58: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Sample/req
      -- 
    if_choice_transition_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1624_branch_ack_1, ack => convTransposeA_CP_3826_elements(58)); -- 
    req_4745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(58), ack => WPIPE_Block0_done_1632_inst_req_0); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	65 
    -- CP-element group 59: 	66 
    -- CP-element group 59: 	68 
    -- CP-element group 59: 	69 
    -- CP-element group 59:  members (20) 
      -- CP-element group 59: 	 branch_block_stmt_1261/if_stmt_1624_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1261/if_stmt_1624_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1624_branch_ack_0, ack => convTransposeA_CP_3826_elements(59)); -- 
    rr_4789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(59), ack => type_cast_1427_inst_req_0); -- 
    cr_4794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(59), ack => type_cast_1427_inst_req_1); -- 
    rr_4812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(59), ack => type_cast_1434_inst_req_0); -- 
    cr_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(59), ack => type_cast_1434_inst_req_1); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Update/req
      -- 
    ack_4746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1632_inst_ack_0, ack => convTransposeA_CP_3826_elements(60)); -- 
    req_4750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(60), ack => WPIPE_Block0_done_1632_inst_req_1); -- 
    -- CP-element group 61:  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (16) 
      -- CP-element group 61: 	 branch_block_stmt_1261/return__
      -- CP-element group 61: 	 branch_block_stmt_1261/branch_block_stmt_1261__exit__
      -- CP-element group 61: 	 branch_block_stmt_1261/assign_stmt_1634__exit__
      -- CP-element group 61: 	 branch_block_stmt_1261/$exit
      -- CP-element group 61: 	 $exit
      -- CP-element group 61: 	 branch_block_stmt_1261/merge_stmt_1636__exit__
      -- CP-element group 61: 	 branch_block_stmt_1261/return___PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_1261/return___PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_1261/merge_stmt_1636_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_1261/merge_stmt_1636_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_1261/merge_stmt_1636_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_1261/merge_stmt_1636_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_1261/assign_stmt_1634/$exit
      -- CP-element group 61: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1261/assign_stmt_1634/WPIPE_Block0_done_1632_Update/ack
      -- 
    ack_4751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1632_inst_ack_1, ack => convTransposeA_CP_3826_elements(61)); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	29 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/$exit
      -- CP-element group 62: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1425_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_req
      -- 
    phi_stmt_1421_req_4762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1421_req_4762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(62), ack => phi_stmt_1421_req_0); -- 
    -- Element group convTransposeA_CP_3826_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => convTransposeA_CP_3826_elements(29), ack => convTransposeA_CP_3826_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  output  delay-element  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	29 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/$exit
      -- CP-element group 63: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1432_konst_delay_trans
      -- CP-element group 63: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_req
      -- 
    phi_stmt_1428_req_4770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1428_req_4770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(63), ack => phi_stmt_1428_req_0); -- 
    -- Element group convTransposeA_CP_3826_elements(63) is a control-delay.
    cp_element_63_delay: control_delay_element  generic map(name => " 63_delay", delay_value => 1)  port map(req => convTransposeA_CP_3826_elements(29), ack => convTransposeA_CP_3826_elements(63), clk => clk, reset =>reset);
    -- CP-element group 64:  join  transition  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	72 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1261/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(62) & convTransposeA_CP_3826_elements(63);
      gj_convTransposeA_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	59 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Sample/ra
      -- 
    ra_4790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_0, ack => convTransposeA_CP_3826_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	59 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/Update/ca
      -- 
    ca_4795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_1, ack => convTransposeA_CP_3826_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/$exit
      -- CP-element group 67: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/$exit
      -- CP-element group 67: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_sources/type_cast_1427/SplitProtocol/$exit
      -- CP-element group 67: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1421/phi_stmt_1421_req
      -- 
    phi_stmt_1421_req_4796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1421_req_4796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(67), ack => phi_stmt_1421_req_1); -- 
    convTransposeA_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(65) & convTransposeA_CP_3826_elements(66);
      gj_convTransposeA_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	59 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Sample/ra
      -- 
    ra_4813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1434_inst_ack_0, ack => convTransposeA_CP_3826_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	59 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/Update/ca
      -- 
    ca_4818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1434_inst_ack_1, ack => convTransposeA_CP_3826_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/$exit
      -- CP-element group 70: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/$exit
      -- CP-element group 70: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_sources/type_cast_1434/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1428/phi_stmt_1428_req
      -- 
    phi_stmt_1428_req_4819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1428_req_4819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(70), ack => phi_stmt_1428_req_1); -- 
    convTransposeA_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(68) & convTransposeA_CP_3826_elements(69);
      gj_convTransposeA_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1261/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(67) & convTransposeA_CP_3826_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  merge  fork  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	64 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1261/merge_stmt_1420_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1261/merge_stmt_1420_PhiAck/$entry
      -- 
    convTransposeA_CP_3826_elements(72) <= OrReduce(convTransposeA_CP_3826_elements(64) & convTransposeA_CP_3826_elements(71));
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1261/merge_stmt_1420_PhiAck/phi_stmt_1421_ack
      -- 
    phi_stmt_1421_ack_4824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1421_ack_0, ack => convTransposeA_CP_3826_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1261/merge_stmt_1420_PhiAck/phi_stmt_1428_ack
      -- 
    phi_stmt_1428_ack_4825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1428_ack_0, ack => convTransposeA_CP_3826_elements(74)); -- 
    -- CP-element group 75:  join  transition  place  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (10) 
      -- CP-element group 75: 	 branch_block_stmt_1261/merge_stmt_1420__exit__
      -- CP-element group 75: 	 branch_block_stmt_1261/assign_stmt_1440_to_assign_stmt_1485__exit__
      -- CP-element group 75: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 75: 	 branch_block_stmt_1261/assign_stmt_1440_to_assign_stmt_1485__entry__
      -- CP-element group 75: 	 branch_block_stmt_1261/assign_stmt_1440_to_assign_stmt_1485/$entry
      -- CP-element group 75: 	 branch_block_stmt_1261/assign_stmt_1440_to_assign_stmt_1485/$exit
      -- CP-element group 75: 	 branch_block_stmt_1261/merge_stmt_1420_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/$entry
      -- CP-element group 75: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/$entry
      -- 
    convTransposeA_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(73) & convTransposeA_CP_3826_elements(74);
      gj_convTransposeA_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	50 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Sample/ra
      -- 
    ra_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1494_inst_ack_0, ack => convTransposeA_CP_3826_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	50 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/Update/ca
      -- 
    ca_4850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1494_inst_ack_1, ack => convTransposeA_CP_3826_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/$exit
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/$exit
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1494/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1261/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_req
      -- 
    phi_stmt_1488_req_4851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1488_req_4851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(78), ack => phi_stmt_1488_req_1); -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3826_elements(76) & convTransposeA_CP_3826_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3826_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/$exit
      -- CP-element group 79: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_sources/type_cast_1492_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1261/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1488/phi_stmt_1488_req
      -- 
    phi_stmt_1488_req_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1488_req_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(79), ack => phi_stmt_1488_req_0); -- 
    -- Element group convTransposeA_CP_3826_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3826_elements(75), ack => convTransposeA_CP_3826_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  merge  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1261/merge_stmt_1487_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1261/merge_stmt_1487_PhiAck/$entry
      -- 
    convTransposeA_CP_3826_elements(80) <= OrReduce(convTransposeA_CP_3826_elements(78) & convTransposeA_CP_3826_elements(79));
    -- CP-element group 81:  fork  transition  place  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	30 
    -- CP-element group 81: 	31 
    -- CP-element group 81: 	33 
    -- CP-element group 81: 	35 
    -- CP-element group 81: 	37 
    -- CP-element group 81: 	38 
    -- CP-element group 81: 	39 
    -- CP-element group 81: 	41 
    -- CP-element group 81: 	43 
    -- CP-element group 81: 	46 
    -- CP-element group 81: 	47 
    -- CP-element group 81: 	48 
    -- CP-element group 81:  members (45) 
      -- CP-element group 81: 	 branch_block_stmt_1261/merge_stmt_1487__exit__
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568__entry__
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1514_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_update_start
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1526_final_index_sum_regn_Update/req
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1527_complete/req
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1531_Update/word_access_complete/word_0/cr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1535_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_update_start
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/array_obj_ref_1547_final_index_sum_regn_Update/req
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/addr_of_1548_complete/req
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/ptr_deref_1551_Update/word_access_complete/word_0/cr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1261/assign_stmt_1501_to_assign_stmt_1568/type_cast_1556_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1261/merge_stmt_1487_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_1261/merge_stmt_1487_PhiAck/phi_stmt_1488_ack
      -- 
    phi_stmt_1488_ack_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1488_ack_0, ack => convTransposeA_CP_3826_elements(81)); -- 
    rr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1514_inst_req_0); -- 
    cr_4427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1514_inst_req_1); -- 
    req_4458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => array_obj_ref_1526_index_offset_req_1); -- 
    req_4473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => addr_of_1527_final_reg_req_1); -- 
    cr_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => ptr_deref_1531_load_0_req_1); -- 
    rr_4532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1535_inst_req_0); -- 
    cr_4537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1535_inst_req_1); -- 
    req_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => array_obj_ref_1547_index_offset_req_1); -- 
    req_4583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => addr_of_1548_final_reg_req_1); -- 
    cr_4633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => ptr_deref_1551_store_0_req_1); -- 
    rr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1556_inst_req_0); -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3826_elements(81), ack => type_cast_1556_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_1313_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1313_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr100_1525_resized : std_logic_vector(13 downto 0);
    signal R_shr100_1525_scaled : std_logic_vector(13 downto 0);
    signal R_shr57102_1546_resized : std_logic_vector(13 downto 0);
    signal R_shr57102_1546_scaled : std_logic_vector(13 downto 0);
    signal add10_1506 : std_logic_vector(15 downto 0);
    signal add50_1511 : std_logic_vector(15 downto 0);
    signal add63_1563 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1526_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1526_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1526_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1526_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1526_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1526_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1547_root_address : std_logic_vector(13 downto 0);
    signal arrayidx59_1549 : std_logic_vector(31 downto 0);
    signal arrayidx_1528 : std_logic_vector(31 downto 0);
    signal call_1264 : std_logic_vector(15 downto 0);
    signal cmp76_1598 : std_logic_vector(0 downto 0);
    signal cmp86_1623 : std_logic_vector(0 downto 0);
    signal cmp_1568 : std_logic_vector(0 downto 0);
    signal conv53_1515 : std_logic_vector(63 downto 0);
    signal conv56_1536 : std_logic_vector(63 downto 0);
    signal conv62_1557 : std_logic_vector(31 downto 0);
    signal conv65_1364 : std_logic_vector(31 downto 0);
    signal conv73_1593 : std_logic_vector(31 downto 0);
    signal conv75_1368 : std_logic_vector(31 downto 0);
    signal conv82_1618 : std_logic_vector(31 downto 0);
    signal conv84_1390 : std_logic_vector(31 downto 0);
    signal div85_1396 : std_logic_vector(31 downto 0);
    signal div_1374 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1382 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1273 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1285 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1295 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1307 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1320 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1332 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1344 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1356 : std_logic_vector(31 downto 0);
    signal inc80_1602 : std_logic_vector(15 downto 0);
    signal inc80x_xinput_dim0x_x2_1607 : std_logic_vector(15 downto 0);
    signal inc_1589 : std_logic_vector(15 downto 0);
    signal indvar_1488 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1581 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1428 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1421 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1614 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1501 : std_logic_vector(15 downto 0);
    signal ptr_deref_1276_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1276_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1276_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1276_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1276_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1288_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1288_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1288_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1288_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1288_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1298_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1298_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1298_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1298_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1298_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1310_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1310_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1310_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1310_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1310_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1323_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1323_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1323_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1323_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1323_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1335_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1335_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1335_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1335_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1335_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1347_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1347_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1347_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1347_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1347_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1359_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1359_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1385_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1385_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1385_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1385_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1385_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1531_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1531_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1531_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1531_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1531_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1551_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1551_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr100_1521 : std_logic_vector(63 downto 0);
    signal shr57102_1542 : std_logic_vector(63 downto 0);
    signal tmp10_1475 : std_logic_vector(15 downto 0);
    signal tmp115_1440 : std_logic_vector(15 downto 0);
    signal tmp116_1445 : std_logic_vector(15 downto 0);
    signal tmp117_1450 : std_logic_vector(15 downto 0);
    signal tmp11_1480 : std_logic_vector(15 downto 0);
    signal tmp12_1485 : std_logic_vector(15 downto 0);
    signal tmp14_1299 : std_logic_vector(15 downto 0);
    signal tmp17_1311 : std_logic_vector(15 downto 0);
    signal tmp1_1277 : std_logic_vector(15 downto 0);
    signal tmp20_1314 : std_logic_vector(15 downto 0);
    signal tmp26_1324 : std_logic_vector(15 downto 0);
    signal tmp29_1336 : std_logic_vector(15 downto 0);
    signal tmp2_1407 : std_logic_vector(15 downto 0);
    signal tmp39_1348 : std_logic_vector(15 downto 0);
    signal tmp3_1455 : std_logic_vector(15 downto 0);
    signal tmp43_1360 : std_logic_vector(15 downto 0);
    signal tmp4_1460 : std_logic_vector(15 downto 0);
    signal tmp54_1532 : std_logic_vector(63 downto 0);
    signal tmp5_1289 : std_logic_vector(15 downto 0);
    signal tmp6_1413 : std_logic_vector(15 downto 0);
    signal tmp7_1418 : std_logic_vector(15 downto 0);
    signal tmp83_1386 : std_logic_vector(15 downto 0);
    signal tmp8_1465 : std_logic_vector(15 downto 0);
    signal tmp9_1470 : std_logic_vector(15 downto 0);
    signal tmp_1402 : std_logic_vector(15 downto 0);
    signal type_cast_1372_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1411_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1425_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1427_wire : std_logic_vector(15 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1434_wire : std_logic_vector(15 downto 0);
    signal type_cast_1492_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1494_wire : std_logic_vector(15 downto 0);
    signal type_cast_1499_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1540_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1561_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1579_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1587_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_1313_word_address_0 <= "0";
    array_obj_ref_1526_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1526_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1526_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1526_resized_base_address <= "00000000000000";
    array_obj_ref_1547_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1547_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1547_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1547_resized_base_address <= "00000000000000";
    iNsTr_10_1382 <= "00000000000000000000000000000011";
    iNsTr_2_1273 <= "00000000000000000000000000000101";
    iNsTr_3_1285 <= "00000000000000000000000000000100";
    iNsTr_4_1295 <= "00000000000000000000000000000000";
    iNsTr_5_1307 <= "00000000000000000000000000000100";
    iNsTr_6_1320 <= "00000000000000000000000000000001";
    iNsTr_7_1332 <= "00000000000000000000000000000101";
    iNsTr_8_1344 <= "00000000000000000000000000000101";
    iNsTr_9_1356 <= "00000000000000000000000000000100";
    ptr_deref_1276_word_offset_0 <= "0000000";
    ptr_deref_1288_word_offset_0 <= "0000000";
    ptr_deref_1298_word_offset_0 <= "0";
    ptr_deref_1310_word_offset_0 <= "0000000";
    ptr_deref_1323_word_offset_0 <= "0";
    ptr_deref_1335_word_offset_0 <= "0000000";
    ptr_deref_1347_word_offset_0 <= "0000000";
    ptr_deref_1359_word_offset_0 <= "0000000";
    ptr_deref_1385_word_offset_0 <= "0000000";
    ptr_deref_1531_word_offset_0 <= "00000000000000";
    ptr_deref_1551_word_offset_0 <= "00000000000000";
    type_cast_1372_wire_constant <= "00000000000000000000000000000001";
    type_cast_1394_wire_constant <= "00000000000000000000000000000001";
    type_cast_1400_wire_constant <= "1111111111111111";
    type_cast_1411_wire_constant <= "1111111111111111";
    type_cast_1425_wire_constant <= "0000000000000000";
    type_cast_1432_wire_constant <= "0000000000000000";
    type_cast_1492_wire_constant <= "0000000000000000";
    type_cast_1499_wire_constant <= "0000000000000100";
    type_cast_1519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1540_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1561_wire_constant <= "00000000000000000000000000000100";
    type_cast_1579_wire_constant <= "0000000000000001";
    type_cast_1587_wire_constant <= "0000000000000001";
    type_cast_1611_wire_constant <= "0000000000000000";
    phi_stmt_1421: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1425_wire_constant & type_cast_1427_wire;
      req <= phi_stmt_1421_req_0 & phi_stmt_1421_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1421",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1421_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1421,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1421
    phi_stmt_1428: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1432_wire_constant & type_cast_1434_wire;
      req <= phi_stmt_1428_req_0 & phi_stmt_1428_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1428",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1428_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1428,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1428
    phi_stmt_1488: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1492_wire_constant & type_cast_1494_wire;
      req <= phi_stmt_1488_req_0 & phi_stmt_1488_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1488",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1488_ack_0,
          idata => idata,
          odata => indvar_1488,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1488
    -- flow-through select operator MUX_1613_inst
    input_dim1x_x2_1614 <= type_cast_1611_wire_constant when (cmp76_1598(0) /=  '0') else inc_1589;
    addr_of_1527_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1527_final_reg_req_0;
      addr_of_1527_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1527_final_reg_req_1;
      addr_of_1527_final_reg_ack_1<= rack(0);
      addr_of_1527_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1527_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1526_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1548_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1548_final_reg_req_0;
      addr_of_1548_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1548_final_reg_req_1;
      addr_of_1548_final_reg_ack_1<= rack(0);
      addr_of_1548_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1548_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1547_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx59_1549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1363_inst_req_0;
      type_cast_1363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1363_inst_req_1;
      type_cast_1363_inst_ack_1<= rack(0);
      type_cast_1363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1367_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1367_inst_req_0;
      type_cast_1367_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1367_inst_req_1;
      type_cast_1367_inst_ack_1<= rack(0);
      type_cast_1367_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1367_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_1289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1368,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1389_inst_req_0;
      type_cast_1389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1389_inst_req_1;
      type_cast_1389_inst_ack_1<= rack(0);
      type_cast_1389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp83_1386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_1390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1427_inst_req_0;
      type_cast_1427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1427_inst_req_1;
      type_cast_1427_inst_ack_1<= rack(0);
      type_cast_1427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1427_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1434_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1434_inst_req_0;
      type_cast_1434_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1434_inst_req_1;
      type_cast_1434_inst_ack_1<= rack(0);
      type_cast_1434_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1434_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc80x_xinput_dim0x_x2_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1434_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1494_inst_req_0;
      type_cast_1494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1494_inst_req_1;
      type_cast_1494_inst_ack_1<= rack(0);
      type_cast_1494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1494_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1514_inst_req_0;
      type_cast_1514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1514_inst_req_1;
      type_cast_1514_inst_ack_1<= rack(0);
      type_cast_1514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add10_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1535_inst_req_0;
      type_cast_1535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1535_inst_req_1;
      type_cast_1535_inst_ack_1<= rack(0);
      type_cast_1535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add50_1511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1556_inst_req_0;
      type_cast_1556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1556_inst_req_1;
      type_cast_1556_inst_ack_1<= rack(0);
      type_cast_1556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1592_inst_req_0;
      type_cast_1592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1592_inst_req_1;
      type_cast_1592_inst_ack_1<= rack(0);
      type_cast_1592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1601_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1601_inst_req_0;
      type_cast_1601_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1601_inst_req_1;
      type_cast_1601_inst_ack_1<= rack(0);
      type_cast_1601_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1601_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp76_1598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc80_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1617_inst_req_0;
      type_cast_1617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1617_inst_req_1;
      type_cast_1617_inst_ack_1<= rack(0);
      type_cast_1617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc80x_xinput_dim0x_x2_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1313_gather_scatter
    process(LOAD_padding_1313_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1313_data_0;
      ov(15 downto 0) := iv;
      tmp20_1314 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1526_index_1_rename
    process(R_shr100_1525_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr100_1525_resized;
      ov(13 downto 0) := iv;
      R_shr100_1525_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1526_index_1_resize
    process(shr100_1521) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr100_1521;
      ov := iv(13 downto 0);
      R_shr100_1525_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1526_root_address_inst
    process(array_obj_ref_1526_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1526_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1526_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_index_1_rename
    process(R_shr57102_1546_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr57102_1546_resized;
      ov(13 downto 0) := iv;
      R_shr57102_1546_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_index_1_resize
    process(shr57102_1542) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr57102_1542;
      ov := iv(13 downto 0);
      R_shr57102_1546_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1547_root_address_inst
    process(array_obj_ref_1547_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1547_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1547_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1276_addr_0
    process(ptr_deref_1276_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1276_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1276_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1276_base_resize
    process(iNsTr_2_1273) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1273;
      ov := iv(6 downto 0);
      ptr_deref_1276_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1276_gather_scatter
    process(ptr_deref_1276_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1276_data_0;
      ov(15 downto 0) := iv;
      tmp1_1277 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1276_root_address_inst
    process(ptr_deref_1276_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1276_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1276_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1288_addr_0
    process(ptr_deref_1288_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1288_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1288_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1288_base_resize
    process(iNsTr_3_1285) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1285;
      ov := iv(6 downto 0);
      ptr_deref_1288_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1288_gather_scatter
    process(ptr_deref_1288_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1288_data_0;
      ov(15 downto 0) := iv;
      tmp5_1289 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1288_root_address_inst
    process(ptr_deref_1288_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1288_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1288_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1298_addr_0
    process(ptr_deref_1298_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1298_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1298_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1298_base_resize
    process(iNsTr_4_1295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1295;
      ov := iv(0 downto 0);
      ptr_deref_1298_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1298_gather_scatter
    process(ptr_deref_1298_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1298_data_0;
      ov(15 downto 0) := iv;
      tmp14_1299 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1298_root_address_inst
    process(ptr_deref_1298_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1298_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1298_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1310_addr_0
    process(ptr_deref_1310_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1310_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1310_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1310_base_resize
    process(iNsTr_5_1307) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1307;
      ov := iv(6 downto 0);
      ptr_deref_1310_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1310_gather_scatter
    process(ptr_deref_1310_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1310_data_0;
      ov(15 downto 0) := iv;
      tmp17_1311 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1310_root_address_inst
    process(ptr_deref_1310_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1310_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1310_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1323_addr_0
    process(ptr_deref_1323_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1323_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1323_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1323_base_resize
    process(iNsTr_6_1320) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1320;
      ov := iv(0 downto 0);
      ptr_deref_1323_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1323_gather_scatter
    process(ptr_deref_1323_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1323_data_0;
      ov(15 downto 0) := iv;
      tmp26_1324 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1323_root_address_inst
    process(ptr_deref_1323_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1323_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1323_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1335_addr_0
    process(ptr_deref_1335_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1335_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1335_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1335_base_resize
    process(iNsTr_7_1332) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1332;
      ov := iv(6 downto 0);
      ptr_deref_1335_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1335_gather_scatter
    process(ptr_deref_1335_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1335_data_0;
      ov(15 downto 0) := iv;
      tmp29_1336 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1335_root_address_inst
    process(ptr_deref_1335_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1335_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1335_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1347_addr_0
    process(ptr_deref_1347_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1347_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1347_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1347_base_resize
    process(iNsTr_8_1344) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1344;
      ov := iv(6 downto 0);
      ptr_deref_1347_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1347_gather_scatter
    process(ptr_deref_1347_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1347_data_0;
      ov(15 downto 0) := iv;
      tmp39_1348 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1347_root_address_inst
    process(ptr_deref_1347_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1347_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1347_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_addr_0
    process(ptr_deref_1359_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1359_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_base_resize
    process(iNsTr_9_1356) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1356;
      ov := iv(6 downto 0);
      ptr_deref_1359_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_gather_scatter
    process(ptr_deref_1359_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_data_0;
      ov(15 downto 0) := iv;
      tmp43_1360 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1359_root_address_inst
    process(ptr_deref_1359_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1359_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1359_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1385_addr_0
    process(ptr_deref_1385_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1385_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1385_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1385_base_resize
    process(iNsTr_10_1382) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1382;
      ov := iv(6 downto 0);
      ptr_deref_1385_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1385_gather_scatter
    process(ptr_deref_1385_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1385_data_0;
      ov(15 downto 0) := iv;
      tmp83_1386 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1385_root_address_inst
    process(ptr_deref_1385_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1385_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1385_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1531_addr_0
    process(ptr_deref_1531_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1531_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1531_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1531_base_resize
    process(arrayidx_1528) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1528;
      ov := iv(13 downto 0);
      ptr_deref_1531_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1531_gather_scatter
    process(ptr_deref_1531_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1531_data_0;
      ov(63 downto 0) := iv;
      tmp54_1532 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1531_root_address_inst
    process(ptr_deref_1531_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1531_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1531_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_addr_0
    process(ptr_deref_1551_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_base_resize
    process(arrayidx59_1549) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx59_1549;
      ov := iv(13 downto 0);
      ptr_deref_1551_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_gather_scatter
    process(tmp54_1532) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp54_1532;
      ov(63 downto 0) := iv;
      ptr_deref_1551_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1551_root_address_inst
    process(ptr_deref_1551_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1551_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1551_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1569_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1568;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1569_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1569_branch_req_0,
          ack0 => if_stmt_1569_branch_ack_0,
          ack1 => if_stmt_1569_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1624_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp86_1623;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1624_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1624_branch_req_0,
          ack0 => if_stmt_1624_branch_ack_0,
          ack1 => if_stmt_1624_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1401_inst
    process(tmp29_1336) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp29_1336, type_cast_1400_wire_constant, tmp_var);
      tmp_1402 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1412_inst
    process(tmp17_1311) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp17_1311, type_cast_1411_wire_constant, tmp_var);
      tmp6_1413 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1444_inst
    process(input_dim1x_x1x_xph_1421, tmp115_1440) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1421, tmp115_1440, tmp_var);
      tmp116_1445 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1459_inst
    process(tmp2_1407, tmp3_1455) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_1407, tmp3_1455, tmp_var);
      tmp4_1460 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1469_inst
    process(tmp7_1418, tmp8_1465) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_1418, tmp8_1465, tmp_var);
      tmp9_1470 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1479_inst
    process(tmp4_1460, tmp10_1475) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_1460, tmp10_1475, tmp_var);
      tmp11_1480 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1505_inst
    process(tmp117_1450, input_dim2x_x1_1501) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp117_1450, input_dim2x_x1_1501, tmp_var);
      add10_1506 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1510_inst
    process(tmp12_1485, input_dim2x_x1_1501) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp12_1485, input_dim2x_x1_1501, tmp_var);
      add50_1511 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1580_inst
    process(indvar_1488) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1488, type_cast_1579_wire_constant, tmp_var);
      indvarx_xnext_1581 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1588_inst
    process(input_dim1x_x1x_xph_1421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1421, type_cast_1587_wire_constant, tmp_var);
      inc_1589 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1606_inst
    process(inc80_1602, input_dim0x_x2x_xph_1428) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc80_1602, input_dim0x_x2x_xph_1428, tmp_var);
      inc80x_xinput_dim0x_x2_1607 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1562_inst
    process(conv62_1557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv62_1557, type_cast_1561_wire_constant, tmp_var);
      add63_1563 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1597_inst
    process(conv73_1593, div_1374) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv73_1593, div_1374, tmp_var);
      cmp76_1598 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1622_inst
    process(conv82_1618, div85_1396) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv82_1618, div85_1396, tmp_var);
      cmp86_1623 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1373_inst
    process(conv75_1368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv75_1368, type_cast_1372_wire_constant, tmp_var);
      div_1374 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1395_inst
    process(conv84_1390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv84_1390, type_cast_1394_wire_constant, tmp_var);
      div85_1396 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1520_inst
    process(conv53_1515) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv53_1515, type_cast_1519_wire_constant, tmp_var);
      shr100_1521 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1541_inst
    process(conv56_1536) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv56_1536, type_cast_1540_wire_constant, tmp_var);
      shr57102_1542 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1439_inst
    process(tmp5_1289, input_dim0x_x2x_xph_1428) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_1289, input_dim0x_x2x_xph_1428, tmp_var);
      tmp115_1440 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1449_inst
    process(tmp1_1277, tmp116_1445) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1277, tmp116_1445, tmp_var);
      tmp117_1450 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1454_inst
    process(tmp26_1324, input_dim1x_x1x_xph_1421) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_1324, input_dim1x_x1x_xph_1421, tmp_var);
      tmp3_1455 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1464_inst
    process(tmp14_1299, input_dim0x_x2x_xph_1428) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1299, input_dim0x_x2x_xph_1428, tmp_var);
      tmp8_1465 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1474_inst
    process(tmp43_1360, tmp9_1470) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp43_1360, tmp9_1470, tmp_var);
      tmp10_1475 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1484_inst
    process(tmp39_1348, tmp11_1480) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp39_1348, tmp11_1480, tmp_var);
      tmp12_1485 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1500_inst
    process(indvar_1488) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1488, type_cast_1499_wire_constant, tmp_var);
      input_dim2x_x1_1501 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1406_inst
    process(tmp_1402, tmp20_1314) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1402, tmp20_1314, tmp_var);
      tmp2_1407 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1417_inst
    process(tmp6_1413, tmp20_1314) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp6_1413, tmp20_1314, tmp_var);
      tmp7_1418 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1567_inst
    process(add63_1563, conv65_1364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add63_1563, conv65_1364, tmp_var);
      cmp_1568 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1526_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr100_1525_scaled;
      array_obj_ref_1526_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1526_index_offset_req_0;
      array_obj_ref_1526_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1526_index_offset_req_1;
      array_obj_ref_1526_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1547_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr57102_1546_scaled;
      array_obj_ref_1547_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1547_index_offset_req_0;
      array_obj_ref_1547_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1547_index_offset_req_1;
      array_obj_ref_1547_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : LOAD_padding_1313_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1313_load_0_req_0;
      LOAD_padding_1313_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1313_load_0_req_1;
      LOAD_padding_1313_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1313_word_address_0;
      LOAD_padding_1313_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1385_load_0 ptr_deref_1288_load_0 ptr_deref_1276_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1385_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1288_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1276_load_0_req_0;
      ptr_deref_1385_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1288_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1276_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1385_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1288_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1276_load_0_req_1;
      ptr_deref_1385_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1288_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1276_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1385_word_address_0 & ptr_deref_1288_word_address_0 & ptr_deref_1276_word_address_0;
      ptr_deref_1385_data_0 <= data_out(47 downto 32);
      ptr_deref_1288_data_0 <= data_out(31 downto 16);
      ptr_deref_1276_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1323_load_0 ptr_deref_1298_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1323_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1298_load_0_req_0;
      ptr_deref_1323_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1298_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1323_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1298_load_0_req_1;
      ptr_deref_1323_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1298_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1323_word_address_0 & ptr_deref_1298_word_address_0;
      ptr_deref_1323_data_0 <= data_out(31 downto 16);
      ptr_deref_1298_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1335_load_0 ptr_deref_1310_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1335_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1310_load_0_req_0;
      ptr_deref_1335_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1310_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1335_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1310_load_0_req_1;
      ptr_deref_1335_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1310_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1335_word_address_0 & ptr_deref_1310_word_address_0;
      ptr_deref_1335_data_0 <= data_out(31 downto 16);
      ptr_deref_1310_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1359_load_0 ptr_deref_1347_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1359_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1347_load_0_req_0;
      ptr_deref_1359_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1347_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1359_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1347_load_0_req_1;
      ptr_deref_1359_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1347_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1359_word_address_0 & ptr_deref_1347_word_address_0;
      ptr_deref_1359_data_0 <= data_out(31 downto 16);
      ptr_deref_1347_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1531_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1531_load_0_req_0;
      ptr_deref_1531_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1531_load_0_req_1;
      ptr_deref_1531_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1531_word_address_0;
      ptr_deref_1531_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1551_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1551_store_0_req_0;
      ptr_deref_1551_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1551_store_0_req_1;
      ptr_deref_1551_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1551_word_address_0;
      data_in <= ptr_deref_1551_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1263_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1263_inst_req_0;
      RPIPE_Block0_start_1263_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1263_inst_req_1;
      RPIPE_Block0_start_1263_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1264 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1632_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1632_inst_req_0;
      WPIPE_Block0_done_1632_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1632_inst_req_1;
      WPIPE_Block0_done_1632_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1264;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4908_start: Boolean;
  signal convTransposeB_CP_4908_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1642_inst_ack_1 : boolean;
  signal ptr_deref_1673_load_0_req_1 : boolean;
  signal RPIPE_Block1_start_1642_inst_req_1 : boolean;
  signal phi_stmt_1796_req_0 : boolean;
  signal ptr_deref_1673_load_0_ack_1 : boolean;
  signal ptr_deref_1695_load_0_req_0 : boolean;
  signal ptr_deref_1683_load_0_req_1 : boolean;
  signal ptr_deref_1673_load_0_req_0 : boolean;
  signal RPIPE_Block1_start_1642_inst_ack_0 : boolean;
  signal ptr_deref_1673_load_0_ack_0 : boolean;
  signal ptr_deref_1683_load_0_req_0 : boolean;
  signal ptr_deref_1655_load_0_ack_1 : boolean;
  signal ptr_deref_1683_load_0_ack_0 : boolean;
  signal ptr_deref_1655_load_0_req_0 : boolean;
  signal ptr_deref_1655_load_0_ack_0 : boolean;
  signal ptr_deref_1655_load_0_req_1 : boolean;
  signal RPIPE_Block1_start_1642_inst_req_0 : boolean;
  signal ptr_deref_1695_load_0_req_1 : boolean;
  signal ptr_deref_1695_load_0_ack_1 : boolean;
  signal ptr_deref_1683_load_0_ack_1 : boolean;
  signal LOAD_padding_1698_load_0_req_0 : boolean;
  signal LOAD_padding_1698_load_0_ack_0 : boolean;
  signal LOAD_padding_1698_load_0_req_1 : boolean;
  signal LOAD_padding_1698_load_0_ack_1 : boolean;
  signal phi_stmt_1802_req_1 : boolean;
  signal type_cast_1808_inst_ack_1 : boolean;
  signal type_cast_1808_inst_req_1 : boolean;
  signal phi_stmt_1862_ack_0 : boolean;
  signal ptr_deref_1708_load_0_req_0 : boolean;
  signal ptr_deref_1708_load_0_ack_0 : boolean;
  signal ptr_deref_1708_load_0_req_1 : boolean;
  signal ptr_deref_1708_load_0_ack_1 : boolean;
  signal ptr_deref_1695_load_0_ack_0 : boolean;
  signal ptr_deref_1720_load_0_req_0 : boolean;
  signal ptr_deref_1720_load_0_ack_0 : boolean;
  signal ptr_deref_1720_load_0_req_1 : boolean;
  signal ptr_deref_1720_load_0_ack_1 : boolean;
  signal phi_stmt_1802_req_0 : boolean;
  signal phi_stmt_1862_req_0 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal ptr_deref_1732_load_0_req_0 : boolean;
  signal ptr_deref_1732_load_0_ack_0 : boolean;
  signal ptr_deref_1732_load_0_req_1 : boolean;
  signal ptr_deref_1732_load_0_ack_1 : boolean;
  signal ptr_deref_1744_load_0_req_0 : boolean;
  signal phi_stmt_1862_req_1 : boolean;
  signal ptr_deref_1744_load_0_ack_0 : boolean;
  signal ptr_deref_1744_load_0_req_1 : boolean;
  signal type_cast_1868_inst_ack_1 : boolean;
  signal ptr_deref_1744_load_0_ack_1 : boolean;
  signal type_cast_1868_inst_req_1 : boolean;
  signal type_cast_1748_inst_req_0 : boolean;
  signal type_cast_1748_inst_ack_0 : boolean;
  signal type_cast_1748_inst_req_1 : boolean;
  signal type_cast_1748_inst_ack_1 : boolean;
  signal type_cast_1868_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2010_inst_ack_1 : boolean;
  signal WPIPE_Block1_done_2010_inst_req_1 : boolean;
  signal ptr_deref_1760_load_0_req_0 : boolean;
  signal ptr_deref_1760_load_0_ack_0 : boolean;
  signal ptr_deref_1760_load_0_req_1 : boolean;
  signal ptr_deref_1760_load_0_ack_1 : boolean;
  signal WPIPE_Block1_done_2010_inst_ack_0 : boolean;
  signal type_cast_1868_inst_req_0 : boolean;
  signal type_cast_1764_inst_req_0 : boolean;
  signal type_cast_1764_inst_ack_0 : boolean;
  signal type_cast_1764_inst_req_1 : boolean;
  signal type_cast_1764_inst_ack_1 : boolean;
  signal type_cast_1888_inst_req_0 : boolean;
  signal type_cast_1888_inst_ack_0 : boolean;
  signal type_cast_1888_inst_req_1 : boolean;
  signal type_cast_1888_inst_ack_1 : boolean;
  signal array_obj_ref_1900_index_offset_req_0 : boolean;
  signal array_obj_ref_1900_index_offset_ack_0 : boolean;
  signal array_obj_ref_1900_index_offset_req_1 : boolean;
  signal array_obj_ref_1900_index_offset_ack_1 : boolean;
  signal type_cast_1799_inst_ack_1 : boolean;
  signal addr_of_1901_final_reg_req_0 : boolean;
  signal addr_of_1901_final_reg_ack_0 : boolean;
  signal addr_of_1901_final_reg_req_1 : boolean;
  signal addr_of_1901_final_reg_ack_1 : boolean;
  signal ptr_deref_1905_load_0_req_0 : boolean;
  signal ptr_deref_1905_load_0_ack_0 : boolean;
  signal WPIPE_Block1_done_2010_inst_req_0 : boolean;
  signal ptr_deref_1905_load_0_req_1 : boolean;
  signal phi_stmt_1802_ack_0 : boolean;
  signal ptr_deref_1905_load_0_ack_1 : boolean;
  signal phi_stmt_1796_ack_0 : boolean;
  signal type_cast_1909_inst_req_0 : boolean;
  signal type_cast_1909_inst_ack_0 : boolean;
  signal type_cast_1909_inst_req_1 : boolean;
  signal type_cast_1909_inst_ack_1 : boolean;
  signal phi_stmt_1796_req_1 : boolean;
  signal type_cast_1801_inst_ack_1 : boolean;
  signal type_cast_1801_inst_req_1 : boolean;
  signal array_obj_ref_1921_index_offset_req_0 : boolean;
  signal array_obj_ref_1921_index_offset_ack_0 : boolean;
  signal type_cast_1799_inst_req_1 : boolean;
  signal array_obj_ref_1921_index_offset_req_1 : boolean;
  signal array_obj_ref_1921_index_offset_ack_1 : boolean;
  signal addr_of_1922_final_reg_req_0 : boolean;
  signal addr_of_1922_final_reg_ack_0 : boolean;
  signal addr_of_1922_final_reg_req_1 : boolean;
  signal addr_of_1922_final_reg_ack_1 : boolean;
  signal type_cast_1799_inst_ack_0 : boolean;
  signal type_cast_1801_inst_ack_0 : boolean;
  signal type_cast_1801_inst_req_0 : boolean;
  signal type_cast_1799_inst_req_0 : boolean;
  signal ptr_deref_1925_store_0_req_0 : boolean;
  signal ptr_deref_1925_store_0_ack_0 : boolean;
  signal ptr_deref_1925_store_0_req_1 : boolean;
  signal ptr_deref_1925_store_0_ack_1 : boolean;
  signal type_cast_1930_inst_req_0 : boolean;
  signal type_cast_1930_inst_ack_0 : boolean;
  signal type_cast_1930_inst_req_1 : boolean;
  signal type_cast_1930_inst_ack_1 : boolean;
  signal if_stmt_1943_branch_req_0 : boolean;
  signal if_stmt_1943_branch_ack_1 : boolean;
  signal if_stmt_1943_branch_ack_0 : boolean;
  signal type_cast_1995_inst_req_0 : boolean;
  signal type_cast_1995_inst_ack_0 : boolean;
  signal type_cast_1995_inst_req_1 : boolean;
  signal type_cast_1995_inst_ack_1 : boolean;
  signal if_stmt_2002_branch_req_0 : boolean;
  signal if_stmt_2002_branch_ack_1 : boolean;
  signal if_stmt_2002_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4908_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4908_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4908_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4908_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4908: Block -- control-path 
    signal convTransposeB_CP_4908_elements: BooleanArray(77 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4908_elements(0) <= convTransposeB_CP_4908_start;
    convTransposeB_CP_4908_symbol <= convTransposeB_CP_4908_elements(55);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1640/$entry
      -- CP-element group 0: 	 branch_block_stmt_1640/assign_stmt_1643__entry__
      -- CP-element group 0: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1640/assign_stmt_1643/$entry
      -- CP-element group 0: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1640/branch_block_stmt_1640__entry__
      -- 
    rr_4956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(0), ack => RPIPE_Block1_start_1642_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Sample/$exit
      -- 
    ra_4957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1642_inst_ack_0, ack => convTransposeB_CP_4908_elements(1)); -- 
    cr_4961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(1), ack => RPIPE_Block1_start_1642_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (259) 
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1643__exit__
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793__entry__
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1643/RPIPE_Block1_start_1642_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1643/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Update/cr
      -- 
    ca_4962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1642_inst_ack_1, ack => convTransposeB_CP_4908_elements(2)); -- 
    cr_5059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1673_load_0_req_1); -- 
    rr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1695_load_0_req_0); -- 
    cr_5109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1683_load_0_req_1); -- 
    rr_5048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1673_load_0_req_0); -- 
    rr_5098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1683_load_0_req_0); -- 
    rr_4998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1655_load_0_req_0); -- 
    cr_5009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1655_load_0_req_1); -- 
    cr_5159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1695_load_0_req_1); -- 
    rr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => LOAD_padding_1698_load_0_req_0); -- 
    cr_5192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => LOAD_padding_1698_load_0_req_1); -- 
    rr_5231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1708_load_0_req_0); -- 
    cr_5242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1708_load_0_req_1); -- 
    rr_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1720_load_0_req_0); -- 
    cr_5292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1720_load_0_req_1); -- 
    rr_5331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1732_load_0_req_0); -- 
    cr_5342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1732_load_0_req_1); -- 
    rr_5381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1744_load_0_req_0); -- 
    cr_5392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1744_load_0_req_1); -- 
    cr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => type_cast_1748_inst_req_1); -- 
    rr_5445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1760_load_0_req_0); -- 
    cr_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => ptr_deref_1760_load_0_req_1); -- 
    cr_5475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(2), ack => type_cast_1764_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Sample/word_access_start/$exit
      -- 
    ra_4999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1655_load_0_ack_0, ack => convTransposeB_CP_4908_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/ptr_deref_1655_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/ptr_deref_1655_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/ptr_deref_1655_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/ptr_deref_1655_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1655_Update/$exit
      -- 
    ca_5010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1655_load_0_ack_1, ack => convTransposeB_CP_4908_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Sample/word_access_start/$exit
      -- 
    ra_5049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1673_load_0_ack_0, ack => convTransposeB_CP_4908_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/ptr_deref_1673_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/ptr_deref_1673_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/ptr_deref_1673_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1673_Update/ptr_deref_1673_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Sample/rr
      -- 
    ca_5060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1673_load_0_ack_1, ack => convTransposeB_CP_4908_elements(6)); -- 
    rr_5406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(6), ack => type_cast_1748_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_sample_completed_
      -- 
    ra_5099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1683_load_0_ack_0, ack => convTransposeB_CP_4908_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	27 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/ptr_deref_1683_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/ptr_deref_1683_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/ptr_deref_1683_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/ptr_deref_1683_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1683_Update/word_access_complete/word_0/ca
      -- 
    ca_5110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1683_load_0_ack_1, ack => convTransposeB_CP_4908_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Sample/word_access_start/word_0/ra
      -- 
    ra_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1695_load_0_ack_0, ack => convTransposeB_CP_4908_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	27 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/ptr_deref_1695_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/ptr_deref_1695_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/ptr_deref_1695_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1695_Update/ptr_deref_1695_Merge/merge_req
      -- 
    ca_5160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1695_load_0_ack_1, ack => convTransposeB_CP_4908_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Sample/word_access_start/$exit
      -- 
    ra_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1698_load_0_ack_0, ack => convTransposeB_CP_4908_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	27 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/LOAD_padding_1698_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/LOAD_padding_1698_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/LOAD_padding_1698_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/LOAD_padding_1698_Update/LOAD_padding_1698_Merge/merge_ack
      -- 
    ca_5193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1698_load_0_ack_1, ack => convTransposeB_CP_4908_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_sample_completed_
      -- 
    ra_5232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1708_load_0_ack_0, ack => convTransposeB_CP_4908_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/ptr_deref_1708_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/ptr_deref_1708_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/ptr_deref_1708_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1708_Update/ptr_deref_1708_Merge/merge_ack
      -- 
    ca_5243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1708_load_0_ack_1, ack => convTransposeB_CP_4908_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Sample/word_access_start/word_0/ra
      -- 
    ra_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_load_0_ack_0, ack => convTransposeB_CP_4908_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	27 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/ptr_deref_1720_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/ptr_deref_1720_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/ptr_deref_1720_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1720_Update/ptr_deref_1720_Merge/merge_ack
      -- 
    ca_5293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_load_0_ack_1, ack => convTransposeB_CP_4908_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Sample/word_access_start/word_0/ra
      -- 
    ra_5332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1732_load_0_ack_0, ack => convTransposeB_CP_4908_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	27 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/ptr_deref_1732_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/ptr_deref_1732_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/ptr_deref_1732_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1732_Update/ptr_deref_1732_Merge/merge_ack
      -- 
    ca_5343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1732_load_0_ack_1, ack => convTransposeB_CP_4908_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Sample/word_access_start/word_0/ra
      -- 
    ra_5382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1744_load_0_ack_0, ack => convTransposeB_CP_4908_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	27 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/ptr_deref_1744_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/ptr_deref_1744_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/ptr_deref_1744_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1744_Update/ptr_deref_1744_Merge/merge_ack
      -- 
    ca_5393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1744_load_0_ack_1, ack => convTransposeB_CP_4908_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Sample/ra
      -- 
    ra_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_0, ack => convTransposeB_CP_4908_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1748_Update/ca
      -- 
    ca_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_1, ack => convTransposeB_CP_4908_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Sample/word_access_start/word_0/ra
      -- 
    ra_5446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1760_load_0_ack_0, ack => convTransposeB_CP_4908_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/ptr_deref_1760_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/ptr_deref_1760_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/ptr_deref_1760_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/ptr_deref_1760_Update/ptr_deref_1760_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Sample/rr
      -- 
    ca_5457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1760_load_0_ack_1, ack => convTransposeB_CP_4908_elements(24)); -- 
    rr_5470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(24), ack => type_cast_1764_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Sample/ra
      -- 
    ra_5471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_0, ack => convTransposeB_CP_4908_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/type_cast_1764_Update/ca
      -- 
    ca_5476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1764_inst_ack_1, ack => convTransposeB_CP_4908_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  place  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	16 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	20 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	8 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	12 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	56 
    -- CP-element group 27: 	57 
    -- CP-element group 27: 	58 
    -- CP-element group 27:  members (14) 
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter
      -- CP-element group 27: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793/$exit
      -- CP-element group 27: 	 branch_block_stmt_1640/assign_stmt_1652_to_assign_stmt_1793__exit__
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/cr
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/$entry
      -- 
    cr_5823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(27), ack => type_cast_1799_inst_req_1); -- 
    rr_5818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(27), ack => type_cast_1799_inst_req_0); -- 
    convTransposeB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(14) & convTransposeB_CP_4908_elements(16) & convTransposeB_CP_4908_elements(18) & convTransposeB_CP_4908_elements(20) & convTransposeB_CP_4908_elements(22) & convTransposeB_CP_4908_elements(26) & convTransposeB_CP_4908_elements(8) & convTransposeB_CP_4908_elements(10) & convTransposeB_CP_4908_elements(12) & convTransposeB_CP_4908_elements(4);
      gj_convTransposeB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	77 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Sample/ra
      -- 
    ra_5491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_0, ack => convTransposeB_CP_4908_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	77 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (16) 
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Sample/req
      -- 
    ca_5496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_1, ack => convTransposeB_CP_4908_elements(29)); -- 
    req_5521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(29), ack => array_obj_ref_1900_index_offset_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	47 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_sample_complete
      -- CP-element group 30: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Sample/ack
      -- 
    ack_5522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1900_index_offset_ack_0, ack => convTransposeB_CP_4908_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	77 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (11) 
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_offset_calculated
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_request/$entry
      -- CP-element group 31: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_request/req
      -- 
    ack_5527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1900_index_offset_ack_1, ack => convTransposeB_CP_4908_elements(31)); -- 
    req_5536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(31), ack => addr_of_1901_final_reg_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_request/$exit
      -- CP-element group 32: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_request/ack
      -- 
    ack_5537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1901_final_reg_ack_0, ack => convTransposeB_CP_4908_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	77 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (24) 
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_complete/ack
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_word_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_address_resized
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_addr_resize/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_addr_resize/$exit
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_addr_resize/base_resize_req
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_addr_resize/base_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_word_addrgen/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_word_addrgen/$exit
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_word_addrgen/root_register_req
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_word_addrgen/root_register_ack
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/word_0/rr
      -- 
    ack_5542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1901_final_reg_ack_1, ack => convTransposeB_CP_4908_elements(33)); -- 
    rr_5575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(33), ack => ptr_deref_1905_load_0_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Sample/word_access_start/word_0/ra
      -- 
    ra_5576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_0, ack => convTransposeB_CP_4908_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	77 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	42 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/ptr_deref_1905_Merge/$entry
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/ptr_deref_1905_Merge/$exit
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_req
      -- CP-element group 35: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_ack
      -- 
    ca_5587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_1, ack => convTransposeB_CP_4908_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	77 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Sample/ra
      -- 
    ra_5601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_0, ack => convTransposeB_CP_4908_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	77 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Sample/req
      -- 
    ca_5606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_1, ack => convTransposeB_CP_4908_elements(37)); -- 
    req_5631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(37), ack => array_obj_ref_1921_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Sample/ack
      -- 
    ack_5632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1921_index_offset_ack_0, ack => convTransposeB_CP_4908_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	77 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_request/req
      -- 
    ack_5637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1921_index_offset_ack_1, ack => convTransposeB_CP_4908_elements(39)); -- 
    req_5646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(39), ack => addr_of_1922_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_request/ack
      -- 
    ack_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1922_final_reg_ack_0, ack => convTransposeB_CP_4908_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	77 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (19) 
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_word_addrgen/root_register_ack
      -- 
    ack_5652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1922_final_reg_ack_1, ack => convTransposeB_CP_4908_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	35 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/ptr_deref_1925_Split/$entry
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/ptr_deref_1925_Split/$exit
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/ptr_deref_1925_Split/split_req
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/ptr_deref_1925_Split/split_ack
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/word_0/rr
      -- 
    rr_5690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(42), ack => ptr_deref_1925_store_0_req_0); -- 
    convTransposeB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(35) & convTransposeB_CP_4908_elements(41);
      gj_convTransposeB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Sample/word_access_start/word_0/ra
      -- 
    ra_5691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1925_store_0_ack_0, ack => convTransposeB_CP_4908_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	77 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/word_0/ca
      -- 
    ca_5702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1925_store_0_ack_1, ack => convTransposeB_CP_4908_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	77 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Sample/ra
      -- 
    ra_5711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_0, ack => convTransposeB_CP_4908_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	77 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Update/ca
      -- 
    ca_5716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_1, ack => convTransposeB_CP_4908_elements(46)); -- 
    -- CP-element group 47:  branch  join  transition  place  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	30 
    -- CP-element group 47: 	38 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (10) 
      -- CP-element group 47: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942__exit__
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943__entry__
      -- CP-element group 47: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/$exit
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_1640/R_cmp_1944_place
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_1640/if_stmt_1943_else_link/$entry
      -- 
    branch_req_5724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(47), ack => if_stmt_1943_branch_req_0); -- 
    convTransposeB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(30) & convTransposeB_CP_4908_elements(38) & convTransposeB_CP_4908_elements(44) & convTransposeB_CP_4908_elements(46);
      gj_convTransposeB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48: 	73 
    -- CP-element group 48:  members (24) 
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody
      -- CP-element group 48: 	 branch_block_stmt_1640/assign_stmt_1955__exit__
      -- CP-element group 48: 	 branch_block_stmt_1640/merge_stmt_1949__exit__
      -- CP-element group 48: 	 branch_block_stmt_1640/assign_stmt_1955__entry__
      -- CP-element group 48: 	 branch_block_stmt_1640/merge_stmt_1949_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_1640/merge_stmt_1949_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_1640/merge_stmt_1949_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_1640/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/merge_stmt_1949_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Update/cr
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/if_stmt_1943_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_1640/if_stmt_1943_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_1640/whilex_xbody_ifx_xthen
      -- CP-element group 48: 	 branch_block_stmt_1640/assign_stmt_1955/$entry
      -- CP-element group 48: 	 branch_block_stmt_1640/assign_stmt_1955/$exit
      -- 
    if_choice_transition_5729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1943_branch_ack_1, ack => convTransposeB_CP_4908_elements(48)); -- 
    cr_5904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(48), ack => type_cast_1868_inst_req_1); -- 
    rr_5899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(48), ack => type_cast_1868_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (18) 
      -- CP-element group 49: 	 branch_block_stmt_1640/merge_stmt_1957__exit__
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001__entry__
      -- CP-element group 49: 	 branch_block_stmt_1640/merge_stmt_1957_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_1640/merge_stmt_1957_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_1640/merge_stmt_1957_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_1640/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_1640/merge_stmt_1957_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_1640/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_1640/if_stmt_1943_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_1640/if_stmt_1943_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_1640/whilex_xbody_ifx_xelse
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/$entry
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Update/cr
      -- 
    else_choice_transition_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1943_branch_ack_0, ack => convTransposeB_CP_4908_elements(49)); -- 
    rr_5749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(49), ack => type_cast_1995_inst_req_0); -- 
    cr_5754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(49), ack => type_cast_1995_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Sample/ra
      -- 
    ra_5750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1995_inst_ack_0, ack => convTransposeB_CP_4908_elements(50)); -- 
    -- CP-element group 51:  branch  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001__exit__
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002__entry__
      -- CP-element group 51: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/$exit
      -- CP-element group 51: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1640/assign_stmt_1963_to_assign_stmt_2001/type_cast_1995_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_dead_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_eval_test/$entry
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_eval_test/$exit
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_eval_test/branch_req
      -- CP-element group 51: 	 branch_block_stmt_1640/R_cmp100_2003_place
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_if_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_1640/if_stmt_2002_else_link/$entry
      -- 
    ca_5755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1995_inst_ack_1, ack => convTransposeB_CP_4908_elements(51)); -- 
    branch_req_5763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(51), ack => if_stmt_2002_branch_req_0); -- 
    -- CP-element group 52:  merge  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (15) 
      -- CP-element group 52: 	 branch_block_stmt_1640/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1640/merge_stmt_2008_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_1640/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_1640/merge_stmt_2008__exit__
      -- CP-element group 52: 	 branch_block_stmt_1640/assign_stmt_2012__entry__
      -- CP-element group 52: 	 branch_block_stmt_1640/merge_stmt_2008_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_1640/merge_stmt_2008_PhiAck/dummy
      -- CP-element group 52: 	 branch_block_stmt_1640/merge_stmt_2008_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1640/if_stmt_2002_if_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1640/if_stmt_2002_if_link/if_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1640/ifx_xelse_whilex_xend
      -- CP-element group 52: 	 branch_block_stmt_1640/assign_stmt_2012/$entry
      -- 
    if_choice_transition_5768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2002_branch_ack_1, ack => convTransposeB_CP_4908_elements(52)); -- 
    req_5785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(52), ack => WPIPE_Block1_done_2010_inst_req_0); -- 
    -- CP-element group 53:  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	61 
    -- CP-element group 53: 	62 
    -- CP-element group 53: 	64 
    -- CP-element group 53: 	65 
    -- CP-element group 53:  members (20) 
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/$entry
      -- CP-element group 53: 	 branch_block_stmt_1640/if_stmt_2002_else_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1640/if_stmt_2002_else_link/else_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter
      -- 
    else_choice_transition_5772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2002_branch_ack_0, ack => convTransposeB_CP_4908_elements(53)); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(53), ack => type_cast_1808_inst_req_1); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(53), ack => type_cast_1808_inst_req_0); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(53), ack => type_cast_1801_inst_req_1); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(53), ack => type_cast_1801_inst_req_0); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Update/req
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_sample_completed_
      -- 
    ack_5786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2010_inst_ack_0, ack => convTransposeB_CP_4908_elements(54)); -- 
    req_5790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(54), ack => WPIPE_Block1_done_2010_inst_req_1); -- 
    -- CP-element group 55:  transition  place  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (16) 
      -- CP-element group 55: 	 branch_block_stmt_1640/$exit
      -- CP-element group 55: 	 branch_block_stmt_1640/branch_block_stmt_1640__exit__
      -- CP-element group 55: 	 $exit
      -- CP-element group 55: 	 branch_block_stmt_1640/assign_stmt_2012__exit__
      -- CP-element group 55: 	 branch_block_stmt_1640/return__
      -- CP-element group 55: 	 branch_block_stmt_1640/merge_stmt_2014__exit__
      -- CP-element group 55: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1640/merge_stmt_2014_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_1640/assign_stmt_2012/WPIPE_Block1_done_2010_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1640/merge_stmt_2014_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_1640/merge_stmt_2014_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_1640/merge_stmt_2014_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_1640/return___PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_1640/return___PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_1640/assign_stmt_2012/$exit
      -- 
    ack_5791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2010_inst_ack_1, ack => convTransposeB_CP_4908_elements(55)); -- 
    -- CP-element group 56:  transition  output  delay-element  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	27 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	60 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_req
      -- CP-element group 56: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1806_konst_delay_trans
      -- CP-element group 56: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/$exit
      -- 
    phi_stmt_1802_req_5802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1802_req_5802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(56), ack => phi_stmt_1802_req_0); -- 
    -- Element group convTransposeB_CP_4908_elements(56) is a control-delay.
    cp_element_56_delay: control_delay_element  generic map(name => " 56_delay", delay_value => 1)  port map(req => convTransposeB_CP_4908_elements(27), ack => convTransposeB_CP_4908_elements(56), clk => clk, reset =>reset);
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	27 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/$exit
      -- 
    ra_5819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_0, ack => convTransposeB_CP_4908_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	27 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/$exit
      -- 
    ca_5824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_1, ack => convTransposeB_CP_4908_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_req
      -- CP-element group 59: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/$exit
      -- CP-element group 59: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/$exit
      -- CP-element group 59: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$exit
      -- CP-element group 59: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/$exit
      -- 
    phi_stmt_1796_req_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1796_req_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(59), ack => phi_stmt_1796_req_0); -- 
    convTransposeB_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(57) & convTransposeB_CP_4908_elements(58);
      gj_convTransposeB_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1640/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(56) & convTransposeB_CP_4908_elements(59);
      gj_convTransposeB_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	53 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Sample/$exit
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_0, ack => convTransposeB_CP_4908_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	53 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/Update/$exit
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_1, ack => convTransposeB_CP_4908_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	67 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_req
      -- CP-element group 63: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/phi_stmt_1802_sources/type_cast_1808/$exit
      -- CP-element group 63: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1802/$exit
      -- 
    phi_stmt_1802_req_5851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1802_req_5851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(63), ack => phi_stmt_1802_req_1); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(61) & convTransposeB_CP_4908_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	53 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Sample/ra
      -- CP-element group 64: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Sample/$exit
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_0, ack => convTransposeB_CP_4908_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	53 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Update/ca
      -- CP-element group 65: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/Update/$exit
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_1, ack => convTransposeB_CP_4908_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/$exit
      -- CP-element group 66: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_req
      -- CP-element group 66: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/SplitProtocol/$exit
      -- CP-element group 66: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1801/$exit
      -- CP-element group 66: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$exit
      -- 
    phi_stmt_1796_req_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1796_req_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(66), ack => phi_stmt_1796_req_1); -- 
    convTransposeB_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(64) & convTransposeB_CP_4908_elements(65);
      gj_convTransposeB_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1640/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(63) & convTransposeB_CP_4908_elements(66);
      gj_convTransposeB_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  merge  fork  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	60 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1640/merge_stmt_1795_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1640/merge_stmt_1795_PhiAck/$entry
      -- 
    convTransposeB_CP_4908_elements(68) <= OrReduce(convTransposeB_CP_4908_elements(60) & convTransposeB_CP_4908_elements(67));
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1640/merge_stmt_1795_PhiAck/phi_stmt_1796_ack
      -- 
    phi_stmt_1796_ack_5879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1796_ack_0, ack => convTransposeB_CP_4908_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1640/merge_stmt_1795_PhiAck/phi_stmt_1802_ack
      -- 
    phi_stmt_1802_ack_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1802_ack_0, ack => convTransposeB_CP_4908_elements(70)); -- 
    -- CP-element group 71:  join  transition  place  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (10) 
      -- CP-element group 71: 	 branch_block_stmt_1640/assign_stmt_1814_to_assign_stmt_1859__exit__
      -- CP-element group 71: 	 branch_block_stmt_1640/assign_stmt_1814_to_assign_stmt_1859__entry__
      -- CP-element group 71: 	 branch_block_stmt_1640/merge_stmt_1795__exit__
      -- CP-element group 71: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 71: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/$entry
      -- CP-element group 71: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_1640/assign_stmt_1814_to_assign_stmt_1859/$entry
      -- CP-element group 71: 	 branch_block_stmt_1640/assign_stmt_1814_to_assign_stmt_1859/$exit
      -- CP-element group 71: 	 branch_block_stmt_1640/merge_stmt_1795_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(69) & convTransposeB_CP_4908_elements(70);
      gj_convTransposeB_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Sample/$exit
      -- 
    ra_5900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1868_inst_ack_0, ack => convTransposeB_CP_4908_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	48 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Update/ca
      -- CP-element group 73: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/Update/$exit
      -- 
    ca_5905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1868_inst_ack_1, ack => convTransposeB_CP_4908_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_req
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1868/$exit
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1862/$exit
      -- CP-element group 74: 	 branch_block_stmt_1640/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1862_req_5906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1862_req_5906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(74), ack => phi_stmt_1862_req_1); -- 
    convTransposeB_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4908_elements(72) & convTransposeB_CP_4908_elements(73);
      gj_convTransposeB_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4908_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_req
      -- CP-element group 75: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/type_cast_1866_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/phi_stmt_1862_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1862/$exit
      -- CP-element group 75: 	 branch_block_stmt_1640/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1862_req_5917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1862_req_5917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(75), ack => phi_stmt_1862_req_0); -- 
    -- Element group convTransposeB_CP_4908_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeB_CP_4908_elements(71), ack => convTransposeB_CP_4908_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  merge  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1640/merge_stmt_1861_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_1640/merge_stmt_1861_PhiReqMerge
      -- 
    convTransposeB_CP_4908_elements(76) <= OrReduce(convTransposeB_CP_4908_elements(74) & convTransposeB_CP_4908_elements(75));
    -- CP-element group 77:  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	28 
    -- CP-element group 77: 	29 
    -- CP-element group 77: 	31 
    -- CP-element group 77: 	33 
    -- CP-element group 77: 	35 
    -- CP-element group 77: 	36 
    -- CP-element group 77: 	37 
    -- CP-element group 77: 	39 
    -- CP-element group 77: 	41 
    -- CP-element group 77: 	44 
    -- CP-element group 77: 	45 
    -- CP-element group 77: 	46 
    -- CP-element group 77:  members (45) 
      -- CP-element group 77: 	 branch_block_stmt_1640/merge_stmt_1861__exit__
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942__entry__
      -- CP-element group 77: 	 branch_block_stmt_1640/merge_stmt_1861_PhiAck/phi_stmt_1862_ack
      -- CP-element group 77: 	 branch_block_stmt_1640/merge_stmt_1861_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1888_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1900_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1901_complete/req
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1905_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1909_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/array_obj_ref_1921_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/addr_of_1922_complete/req
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/ptr_deref_1925_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1640/assign_stmt_1875_to_assign_stmt_1942/type_cast_1930_Update/cr
      -- 
    phi_stmt_1862_ack_5922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1862_ack_0, ack => convTransposeB_CP_4908_elements(77)); -- 
    rr_5490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1888_inst_req_0); -- 
    cr_5495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1888_inst_req_1); -- 
    req_5526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => array_obj_ref_1900_index_offset_req_1); -- 
    req_5541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => addr_of_1901_final_reg_req_1); -- 
    cr_5586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => ptr_deref_1905_load_0_req_1); -- 
    rr_5600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1909_inst_req_0); -- 
    cr_5605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1909_inst_req_1); -- 
    req_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => array_obj_ref_1921_index_offset_req_1); -- 
    req_5651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => addr_of_1922_final_reg_req_1); -- 
    cr_5701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => ptr_deref_1925_store_0_req_1); -- 
    rr_5710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1930_inst_req_0); -- 
    cr_5715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4908_elements(77), ack => type_cast_1930_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_1698_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1698_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr114_1899_resized : std_logic_vector(13 downto 0);
    signal R_shr114_1899_scaled : std_logic_vector(13 downto 0);
    signal R_shr67116_1920_resized : std_logic_vector(13 downto 0);
    signal R_shr67116_1920_scaled : std_logic_vector(13 downto 0);
    signal add20_1880 : std_logic_vector(15 downto 0);
    signal add60_1885 : std_logic_vector(15 downto 0);
    signal add73_1937 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1900_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1900_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1921_root_address : std_logic_vector(13 downto 0);
    signal arrayidx69_1923 : std_logic_vector(31 downto 0);
    signal arrayidx_1902 : std_logic_vector(31 downto 0);
    signal call_1643 : std_logic_vector(15 downto 0);
    signal cmp100_2001 : std_logic_vector(0 downto 0);
    signal cmp86_1968 : std_logic_vector(0 downto 0);
    signal cmp_1942 : std_logic_vector(0 downto 0);
    signal conv63_1889 : std_logic_vector(63 downto 0);
    signal conv66_1910 : std_logic_vector(63 downto 0);
    signal conv72_1931 : std_logic_vector(31 downto 0);
    signal conv75_1749 : std_logic_vector(31 downto 0);
    signal conv96_1996 : std_logic_vector(31 downto 0);
    signal conv98_1765 : std_logic_vector(31 downto 0);
    signal div93_1980 : std_logic_vector(15 downto 0);
    signal div99_1771 : std_logic_vector(31 downto 0);
    signal div_1662 : std_logic_vector(15 downto 0);
    signal iNsTr_10_1757 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1652 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1670 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1680 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1692 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1705 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1717 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1729 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1741 : std_logic_vector(31 downto 0);
    signal inc90_1974 : std_logic_vector(15 downto 0);
    signal inc_1963 : std_logic_vector(15 downto 0);
    signal indvar_1862 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1955 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_1992 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1802 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1796 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1986 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1875 : std_logic_vector(15 downto 0);
    signal ptr_deref_1655_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1655_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1655_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1655_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1655_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1673_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1673_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1673_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1673_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1673_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1683_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1683_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1683_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1683_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1683_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1695_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1695_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1695_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1695_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1695_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1708_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1708_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1708_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1708_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1708_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1720_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1720_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1720_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1720_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1720_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1732_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1732_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1732_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1732_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1732_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1744_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1744_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1744_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1744_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1744_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1760_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1760_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1905_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1905_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1905_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1925_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1925_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1925_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1925_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1925_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1925_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr114_1895 : std_logic_vector(63 downto 0);
    signal shr67116_1916 : std_logic_vector(63 downto 0);
    signal tmp10_1844 : std_logic_vector(15 downto 0);
    signal tmp11_1674 : std_logic_vector(15 downto 0);
    signal tmp12_1849 : std_logic_vector(15 downto 0);
    signal tmp130_1814 : std_logic_vector(15 downto 0);
    signal tmp131_1819 : std_logic_vector(15 downto 0);
    signal tmp132_1824 : std_logic_vector(15 downto 0);
    signal tmp13_1854 : std_logic_vector(15 downto 0);
    signal tmp14_1859 : std_logic_vector(15 downto 0);
    signal tmp24_1684 : std_logic_vector(15 downto 0);
    signal tmp27_1696 : std_logic_vector(15 downto 0);
    signal tmp30_1699 : std_logic_vector(15 downto 0);
    signal tmp36_1709 : std_logic_vector(15 downto 0);
    signal tmp39_1721 : std_logic_vector(15 downto 0);
    signal tmp3_1777 : std_logic_vector(15 downto 0);
    signal tmp49_1733 : std_logic_vector(15 downto 0);
    signal tmp4_1782 : std_logic_vector(15 downto 0);
    signal tmp53_1745 : std_logic_vector(15 downto 0);
    signal tmp5_1829 : std_logic_vector(15 downto 0);
    signal tmp64_1906 : std_logic_vector(63 downto 0);
    signal tmp6_1834 : std_logic_vector(15 downto 0);
    signal tmp7_1788 : std_logic_vector(15 downto 0);
    signal tmp8_1793 : std_logic_vector(15 downto 0);
    signal tmp97_1761 : std_logic_vector(15 downto 0);
    signal tmp9_1839 : std_logic_vector(15 downto 0);
    signal tmp_1656 : std_logic_vector(15 downto 0);
    signal type_cast_1660_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1769_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1775_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1786_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1799_wire : std_logic_vector(15 downto 0);
    signal type_cast_1801_wire : std_logic_vector(15 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1808_wire : std_logic_vector(15 downto 0);
    signal type_cast_1866_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1868_wire : std_logic_vector(15 downto 0);
    signal type_cast_1873_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1893_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1953_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1961_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1972_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1978_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_1698_word_address_0 <= "0";
    array_obj_ref_1900_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1900_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1900_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1900_resized_base_address <= "00000000000000";
    array_obj_ref_1921_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1921_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1921_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1921_resized_base_address <= "00000000000000";
    iNsTr_10_1757 <= "00000000000000000000000000000011";
    iNsTr_2_1652 <= "00000000000000000000000000000100";
    iNsTr_3_1670 <= "00000000000000000000000000000101";
    iNsTr_4_1680 <= "00000000000000000000000000000000";
    iNsTr_5_1692 <= "00000000000000000000000000000100";
    iNsTr_6_1705 <= "00000000000000000000000000000001";
    iNsTr_7_1717 <= "00000000000000000000000000000101";
    iNsTr_8_1729 <= "00000000000000000000000000000101";
    iNsTr_9_1741 <= "00000000000000000000000000000100";
    ptr_deref_1655_word_offset_0 <= "0000000";
    ptr_deref_1673_word_offset_0 <= "0000000";
    ptr_deref_1683_word_offset_0 <= "0";
    ptr_deref_1695_word_offset_0 <= "0000000";
    ptr_deref_1708_word_offset_0 <= "0";
    ptr_deref_1720_word_offset_0 <= "0000000";
    ptr_deref_1732_word_offset_0 <= "0000000";
    ptr_deref_1744_word_offset_0 <= "0000000";
    ptr_deref_1760_word_offset_0 <= "0000000";
    ptr_deref_1905_word_offset_0 <= "00000000000000";
    ptr_deref_1925_word_offset_0 <= "00000000000000";
    type_cast_1660_wire_constant <= "0000000000000001";
    type_cast_1769_wire_constant <= "00000000000000000000000000000001";
    type_cast_1775_wire_constant <= "1111111111111111";
    type_cast_1786_wire_constant <= "1111111111111111";
    type_cast_1806_wire_constant <= "0000000000000000";
    type_cast_1866_wire_constant <= "0000000000000000";
    type_cast_1873_wire_constant <= "0000000000000100";
    type_cast_1893_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1914_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1935_wire_constant <= "00000000000000000000000000000100";
    type_cast_1953_wire_constant <= "0000000000000001";
    type_cast_1961_wire_constant <= "0000000000000001";
    type_cast_1972_wire_constant <= "0000000000000001";
    type_cast_1978_wire_constant <= "0000000000000001";
    phi_stmt_1796: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1799_wire & type_cast_1801_wire;
      req <= phi_stmt_1796_req_0 & phi_stmt_1796_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1796",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1796_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1796,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1796
    phi_stmt_1802: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1806_wire_constant & type_cast_1808_wire;
      req <= phi_stmt_1802_req_0 & phi_stmt_1802_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1802",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1802_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1802,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1802
    phi_stmt_1862: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1866_wire_constant & type_cast_1868_wire;
      req <= phi_stmt_1862_req_0 & phi_stmt_1862_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1862",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1862_ack_0,
          idata => idata,
          odata => indvar_1862,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1862
    -- flow-through select operator MUX_1985_inst
    input_dim1x_x2_1986 <= div93_1980 when (cmp86_1968(0) /=  '0') else inc_1963;
    -- flow-through select operator MUX_1991_inst
    input_dim0x_x0_1992 <= inc90_1974 when (cmp86_1968(0) /=  '0') else input_dim0x_x2x_xph_1802;
    addr_of_1901_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1901_final_reg_req_0;
      addr_of_1901_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1901_final_reg_req_1;
      addr_of_1901_final_reg_ack_1<= rack(0);
      addr_of_1901_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1901_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1900_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1902,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1922_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1922_final_reg_req_0;
      addr_of_1922_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1922_final_reg_req_1;
      addr_of_1922_final_reg_ack_1<= rack(0);
      addr_of_1922_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1922_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1921_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx69_1923,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1748_inst_req_0;
      type_cast_1748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1748_inst_req_1;
      type_cast_1748_inst_ack_1<= rack(0);
      type_cast_1748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_1674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1764_inst_req_0;
      type_cast_1764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1764_inst_req_1;
      type_cast_1764_inst_ack_1<= rack(0);
      type_cast_1764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp97_1761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_1765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1799_inst_req_0;
      type_cast_1799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1799_inst_req_1;
      type_cast_1799_inst_ack_1<= rack(0);
      type_cast_1799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1801_inst_req_0;
      type_cast_1801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1801_inst_req_1;
      type_cast_1801_inst_ack_1<= rack(0);
      type_cast_1801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1986,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1801_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1808_inst_req_0;
      type_cast_1808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1808_inst_req_1;
      type_cast_1808_inst_ack_1<= rack(0);
      type_cast_1808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1992,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1808_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1868_inst_req_0;
      type_cast_1868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1868_inst_req_1;
      type_cast_1868_inst_ack_1<= rack(0);
      type_cast_1868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1955,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1868_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1888_inst_req_0;
      type_cast_1888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1888_inst_req_1;
      type_cast_1888_inst_ack_1<= rack(0);
      type_cast_1888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add20_1880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_1889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1909_inst_req_0;
      type_cast_1909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1909_inst_req_1;
      type_cast_1909_inst_ack_1<= rack(0);
      type_cast_1909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add60_1885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1910,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1930_inst_req_0;
      type_cast_1930_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1930_inst_req_1;
      type_cast_1930_inst_ack_1<= rack(0);
      type_cast_1930_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1930_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1931,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1995_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1995_inst_req_0;
      type_cast_1995_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1995_inst_req_1;
      type_cast_1995_inst_ack_1<= rack(0);
      type_cast_1995_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1995_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1992,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_1996,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1698_gather_scatter
    process(LOAD_padding_1698_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1698_data_0;
      ov(15 downto 0) := iv;
      tmp30_1699 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_index_1_rename
    process(R_shr114_1899_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr114_1899_resized;
      ov(13 downto 0) := iv;
      R_shr114_1899_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_index_1_resize
    process(shr114_1895) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr114_1895;
      ov := iv(13 downto 0);
      R_shr114_1899_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1900_root_address_inst
    process(array_obj_ref_1900_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1900_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1900_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1921_index_1_rename
    process(R_shr67116_1920_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr67116_1920_resized;
      ov(13 downto 0) := iv;
      R_shr67116_1920_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1921_index_1_resize
    process(shr67116_1916) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr67116_1916;
      ov := iv(13 downto 0);
      R_shr67116_1920_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1921_root_address_inst
    process(array_obj_ref_1921_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1921_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1921_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1655_addr_0
    process(ptr_deref_1655_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1655_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1655_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1655_base_resize
    process(iNsTr_2_1652) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1652;
      ov := iv(6 downto 0);
      ptr_deref_1655_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1655_gather_scatter
    process(ptr_deref_1655_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1655_data_0;
      ov(15 downto 0) := iv;
      tmp_1656 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1655_root_address_inst
    process(ptr_deref_1655_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1655_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1655_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_addr_0
    process(ptr_deref_1673_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1673_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1673_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_base_resize
    process(iNsTr_3_1670) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1670;
      ov := iv(6 downto 0);
      ptr_deref_1673_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_gather_scatter
    process(ptr_deref_1673_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1673_data_0;
      ov(15 downto 0) := iv;
      tmp11_1674 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_root_address_inst
    process(ptr_deref_1673_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1673_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1673_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1683_addr_0
    process(ptr_deref_1683_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1683_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1683_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1683_base_resize
    process(iNsTr_4_1680) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1680;
      ov := iv(0 downto 0);
      ptr_deref_1683_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1683_gather_scatter
    process(ptr_deref_1683_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1683_data_0;
      ov(15 downto 0) := iv;
      tmp24_1684 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1683_root_address_inst
    process(ptr_deref_1683_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1683_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1683_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1695_addr_0
    process(ptr_deref_1695_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1695_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1695_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1695_base_resize
    process(iNsTr_5_1692) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1692;
      ov := iv(6 downto 0);
      ptr_deref_1695_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1695_gather_scatter
    process(ptr_deref_1695_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1695_data_0;
      ov(15 downto 0) := iv;
      tmp27_1696 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1695_root_address_inst
    process(ptr_deref_1695_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1695_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1695_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1708_addr_0
    process(ptr_deref_1708_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1708_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1708_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1708_base_resize
    process(iNsTr_6_1705) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1705;
      ov := iv(0 downto 0);
      ptr_deref_1708_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1708_gather_scatter
    process(ptr_deref_1708_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1708_data_0;
      ov(15 downto 0) := iv;
      tmp36_1709 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1708_root_address_inst
    process(ptr_deref_1708_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1708_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1708_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_addr_0
    process(ptr_deref_1720_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1720_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_base_resize
    process(iNsTr_7_1717) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1717;
      ov := iv(6 downto 0);
      ptr_deref_1720_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_gather_scatter
    process(ptr_deref_1720_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_data_0;
      ov(15 downto 0) := iv;
      tmp39_1721 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_root_address_inst
    process(ptr_deref_1720_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1720_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1732_addr_0
    process(ptr_deref_1732_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1732_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1732_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1732_base_resize
    process(iNsTr_8_1729) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1729;
      ov := iv(6 downto 0);
      ptr_deref_1732_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1732_gather_scatter
    process(ptr_deref_1732_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1732_data_0;
      ov(15 downto 0) := iv;
      tmp49_1733 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1732_root_address_inst
    process(ptr_deref_1732_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1732_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1732_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_addr_0
    process(ptr_deref_1744_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1744_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1744_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_base_resize
    process(iNsTr_9_1741) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1741;
      ov := iv(6 downto 0);
      ptr_deref_1744_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_gather_scatter
    process(ptr_deref_1744_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1744_data_0;
      ov(15 downto 0) := iv;
      tmp53_1745 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1744_root_address_inst
    process(ptr_deref_1744_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1744_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1744_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1760_addr_0
    process(ptr_deref_1760_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1760_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1760_base_resize
    process(iNsTr_10_1757) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1757;
      ov := iv(6 downto 0);
      ptr_deref_1760_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1760_gather_scatter
    process(ptr_deref_1760_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_data_0;
      ov(15 downto 0) := iv;
      tmp97_1761 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1760_root_address_inst
    process(ptr_deref_1760_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1760_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1760_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_addr_0
    process(ptr_deref_1905_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1905_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_base_resize
    process(arrayidx_1902) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1902;
      ov := iv(13 downto 0);
      ptr_deref_1905_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_gather_scatter
    process(ptr_deref_1905_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_data_0;
      ov(63 downto 0) := iv;
      tmp64_1906 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_root_address_inst
    process(ptr_deref_1905_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1905_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1925_addr_0
    process(ptr_deref_1925_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1925_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1925_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1925_base_resize
    process(arrayidx69_1923) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx69_1923;
      ov := iv(13 downto 0);
      ptr_deref_1925_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1925_gather_scatter
    process(tmp64_1906) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp64_1906;
      ov(63 downto 0) := iv;
      ptr_deref_1925_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1925_root_address_inst
    process(ptr_deref_1925_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1925_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1925_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1943_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1942;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1943_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1943_branch_req_0,
          ack0 => if_stmt_1943_branch_ack_0,
          ack1 => if_stmt_1943_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2002_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp100_2001;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2002_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2002_branch_req_0,
          ack0 => if_stmt_2002_branch_ack_0,
          ack1 => if_stmt_2002_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1776_inst
    process(tmp39_1721) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp39_1721, type_cast_1775_wire_constant, tmp_var);
      tmp3_1777 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1787_inst
    process(tmp27_1696) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp27_1696, type_cast_1786_wire_constant, tmp_var);
      tmp7_1788 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1818_inst
    process(input_dim1x_x1x_xph_1796, tmp130_1814) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1796, tmp130_1814, tmp_var);
      tmp131_1819 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1833_inst
    process(tmp4_1782, tmp5_1829) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_1782, tmp5_1829, tmp_var);
      tmp6_1834 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1843_inst
    process(tmp8_1793, tmp9_1839) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_1793, tmp9_1839, tmp_var);
      tmp10_1844 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1853_inst
    process(tmp6_1834, tmp12_1849) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_1834, tmp12_1849, tmp_var);
      tmp13_1854 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1879_inst
    process(tmp132_1824, input_dim2x_x1_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp132_1824, input_dim2x_x1_1875, tmp_var);
      add20_1880 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1884_inst
    process(tmp14_1859, input_dim2x_x1_1875) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_1859, input_dim2x_x1_1875, tmp_var);
      add60_1885 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1954_inst
    process(indvar_1862) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1862, type_cast_1953_wire_constant, tmp_var);
      indvarx_xnext_1955 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1962_inst
    process(input_dim1x_x1x_xph_1796) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1796, type_cast_1961_wire_constant, tmp_var);
      inc_1963 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1973_inst
    process(input_dim0x_x2x_xph_1802) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1802, type_cast_1972_wire_constant, tmp_var);
      inc90_1974 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1936_inst
    process(conv72_1931) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv72_1931, type_cast_1935_wire_constant, tmp_var);
      add73_1937 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1967_inst
    process(inc_1963, tmp_1656) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1963, tmp_1656, tmp_var);
      cmp86_1968 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2000_inst
    process(conv96_1996, div99_1771) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv96_1996, div99_1771, tmp_var);
      cmp100_2001 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1661_inst
    process(tmp_1656) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1656, type_cast_1660_wire_constant, tmp_var);
      div_1662 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1979_inst
    process(tmp_1656) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1656, type_cast_1978_wire_constant, tmp_var);
      div93_1980 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1770_inst
    process(conv98_1765) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv98_1765, type_cast_1769_wire_constant, tmp_var);
      div99_1771 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1894_inst
    process(conv63_1889) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv63_1889, type_cast_1893_wire_constant, tmp_var);
      shr114_1895 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1915_inst
    process(conv66_1910) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv66_1910, type_cast_1914_wire_constant, tmp_var);
      shr67116_1916 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1813_inst
    process(tmp_1656, input_dim0x_x2x_xph_1802) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1656, input_dim0x_x2x_xph_1802, tmp_var);
      tmp130_1814 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1823_inst
    process(tmp11_1674, tmp131_1819) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_1674, tmp131_1819, tmp_var);
      tmp132_1824 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1828_inst
    process(tmp36_1709, input_dim1x_x1x_xph_1796) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp36_1709, input_dim1x_x1x_xph_1796, tmp_var);
      tmp5_1829 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1838_inst
    process(tmp24_1684, input_dim0x_x2x_xph_1802) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp24_1684, input_dim0x_x2x_xph_1802, tmp_var);
      tmp9_1839 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1848_inst
    process(tmp53_1745, tmp10_1844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp53_1745, tmp10_1844, tmp_var);
      tmp12_1849 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1858_inst
    process(tmp49_1733, tmp13_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp49_1733, tmp13_1854, tmp_var);
      tmp14_1859 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1874_inst
    process(indvar_1862) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1862, type_cast_1873_wire_constant, tmp_var);
      input_dim2x_x1_1875 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1781_inst
    process(tmp3_1777, tmp30_1699) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_1777, tmp30_1699, tmp_var);
      tmp4_1782 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1792_inst
    process(tmp7_1788, tmp30_1699) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_1788, tmp30_1699, tmp_var);
      tmp8_1793 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1941_inst
    process(add73_1937, conv75_1749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add73_1937, conv75_1749, tmp_var);
      cmp_1942 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_1900_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr114_1899_scaled;
      array_obj_ref_1900_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1900_index_offset_req_0;
      array_obj_ref_1900_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1900_index_offset_req_1;
      array_obj_ref_1900_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_1921_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr67116_1920_scaled;
      array_obj_ref_1921_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1921_index_offset_req_0;
      array_obj_ref_1921_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1921_index_offset_req_1;
      array_obj_ref_1921_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : LOAD_padding_1698_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1698_load_0_req_0;
      LOAD_padding_1698_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1698_load_0_req_1;
      LOAD_padding_1698_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1698_word_address_0;
      LOAD_padding_1698_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1655_load_0 ptr_deref_1760_load_0 ptr_deref_1673_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1655_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1760_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1673_load_0_req_0;
      ptr_deref_1655_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1760_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1673_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1655_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1760_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1673_load_0_req_1;
      ptr_deref_1655_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1760_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1673_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1655_word_address_0 & ptr_deref_1760_word_address_0 & ptr_deref_1673_word_address_0;
      ptr_deref_1655_data_0 <= data_out(47 downto 32);
      ptr_deref_1760_data_0 <= data_out(31 downto 16);
      ptr_deref_1673_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1683_load_0 ptr_deref_1708_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1683_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1708_load_0_req_0;
      ptr_deref_1683_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1708_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1683_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1708_load_0_req_1;
      ptr_deref_1683_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1708_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1683_word_address_0 & ptr_deref_1708_word_address_0;
      ptr_deref_1683_data_0 <= data_out(31 downto 16);
      ptr_deref_1708_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1720_load_0 ptr_deref_1695_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1720_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1695_load_0_req_0;
      ptr_deref_1720_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1695_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1720_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1695_load_0_req_1;
      ptr_deref_1720_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1695_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1720_word_address_0 & ptr_deref_1695_word_address_0;
      ptr_deref_1720_data_0 <= data_out(31 downto 16);
      ptr_deref_1695_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1732_load_0 ptr_deref_1744_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1732_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1744_load_0_req_0;
      ptr_deref_1732_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1744_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1732_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1744_load_0_req_1;
      ptr_deref_1732_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1744_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1732_word_address_0 & ptr_deref_1744_word_address_0;
      ptr_deref_1732_data_0 <= data_out(31 downto 16);
      ptr_deref_1744_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1905_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1905_load_0_req_0;
      ptr_deref_1905_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1905_load_0_req_1;
      ptr_deref_1905_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1905_word_address_0;
      ptr_deref_1905_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1925_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1925_store_0_req_0;
      ptr_deref_1925_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1925_store_0_req_1;
      ptr_deref_1925_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1925_word_address_0;
      data_in <= ptr_deref_1925_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1642_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1642_inst_req_0;
      RPIPE_Block1_start_1642_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1642_inst_req_1;
      RPIPE_Block1_start_1642_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1643 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2010_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2010_inst_req_0;
      WPIPE_Block1_done_2010_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2010_inst_req_1;
      WPIPE_Block1_done_2010_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1643;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5963_start: Boolean;
  signal convTransposeC_CP_5963_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2033_load_0_ack_0 : boolean;
  signal type_cast_2177_inst_ack_0 : boolean;
  signal type_cast_2177_inst_req_0 : boolean;
  signal ptr_deref_2033_load_0_ack_1 : boolean;
  signal ptr_deref_2033_load_0_req_1 : boolean;
  signal RPIPE_Block2_start_2020_inst_ack_1 : boolean;
  signal ptr_deref_2033_load_0_req_0 : boolean;
  signal RPIPE_Block2_start_2020_inst_req_1 : boolean;
  signal ptr_deref_2051_load_0_req_0 : boolean;
  signal ptr_deref_2051_load_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2020_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2020_inst_ack_0 : boolean;
  signal phi_stmt_2240_ack_0 : boolean;
  signal type_cast_2184_inst_req_0 : boolean;
  signal type_cast_2184_inst_ack_0 : boolean;
  signal type_cast_2177_inst_req_1 : boolean;
  signal phi_stmt_2174_ack_0 : boolean;
  signal ptr_deref_2051_load_0_req_1 : boolean;
  signal ptr_deref_2051_load_0_ack_1 : boolean;
  signal ptr_deref_2063_load_0_req_0 : boolean;
  signal ptr_deref_2063_load_0_ack_0 : boolean;
  signal ptr_deref_2063_load_0_req_1 : boolean;
  signal ptr_deref_2063_load_0_ack_1 : boolean;
  signal ptr_deref_2073_load_0_req_0 : boolean;
  signal ptr_deref_2073_load_0_ack_0 : boolean;
  signal ptr_deref_2073_load_0_req_1 : boolean;
  signal ptr_deref_2073_load_0_ack_1 : boolean;
  signal ptr_deref_2085_load_0_req_0 : boolean;
  signal ptr_deref_2085_load_0_ack_0 : boolean;
  signal ptr_deref_2085_load_0_req_1 : boolean;
  signal ptr_deref_2085_load_0_ack_1 : boolean;
  signal LOAD_padding_2088_load_0_req_0 : boolean;
  signal LOAD_padding_2088_load_0_ack_0 : boolean;
  signal LOAD_padding_2088_load_0_req_1 : boolean;
  signal LOAD_padding_2088_load_0_ack_1 : boolean;
  signal ptr_deref_2098_load_0_req_0 : boolean;
  signal ptr_deref_2098_load_0_ack_0 : boolean;
  signal ptr_deref_2098_load_0_req_1 : boolean;
  signal ptr_deref_2098_load_0_ack_1 : boolean;
  signal ptr_deref_2110_load_0_req_0 : boolean;
  signal ptr_deref_2110_load_0_ack_0 : boolean;
  signal ptr_deref_2110_load_0_req_1 : boolean;
  signal ptr_deref_2110_load_0_ack_1 : boolean;
  signal ptr_deref_2122_load_0_req_0 : boolean;
  signal ptr_deref_2122_load_0_ack_0 : boolean;
  signal ptr_deref_2122_load_0_req_1 : boolean;
  signal ptr_deref_2122_load_0_ack_1 : boolean;
  signal ptr_deref_2134_load_0_req_0 : boolean;
  signal ptr_deref_2134_load_0_ack_0 : boolean;
  signal ptr_deref_2134_load_0_req_1 : boolean;
  signal ptr_deref_2134_load_0_ack_1 : boolean;
  signal type_cast_2138_inst_req_0 : boolean;
  signal type_cast_2138_inst_ack_0 : boolean;
  signal type_cast_2138_inst_req_1 : boolean;
  signal type_cast_2138_inst_ack_1 : boolean;
  signal type_cast_2142_inst_req_0 : boolean;
  signal type_cast_2142_inst_ack_0 : boolean;
  signal type_cast_2142_inst_req_1 : boolean;
  signal type_cast_2142_inst_ack_1 : boolean;
  signal phi_stmt_2240_req_1 : boolean;
  signal type_cast_2266_inst_req_0 : boolean;
  signal type_cast_2266_inst_ack_0 : boolean;
  signal type_cast_2266_inst_req_1 : boolean;
  signal type_cast_2266_inst_ack_1 : boolean;
  signal phi_stmt_2181_req_1 : boolean;
  signal array_obj_ref_2278_index_offset_req_0 : boolean;
  signal array_obj_ref_2278_index_offset_ack_0 : boolean;
  signal array_obj_ref_2278_index_offset_req_1 : boolean;
  signal array_obj_ref_2278_index_offset_ack_1 : boolean;
  signal phi_stmt_2240_req_0 : boolean;
  signal addr_of_2279_final_reg_req_0 : boolean;
  signal addr_of_2279_final_reg_ack_0 : boolean;
  signal addr_of_2279_final_reg_req_1 : boolean;
  signal addr_of_2279_final_reg_ack_1 : boolean;
  signal type_cast_2243_inst_ack_1 : boolean;
  signal type_cast_2243_inst_req_1 : boolean;
  signal type_cast_2243_inst_ack_0 : boolean;
  signal type_cast_2243_inst_req_0 : boolean;
  signal type_cast_2186_inst_ack_1 : boolean;
  signal phi_stmt_2181_req_0 : boolean;
  signal type_cast_2184_inst_ack_1 : boolean;
  signal ptr_deref_2283_load_0_req_0 : boolean;
  signal ptr_deref_2283_load_0_ack_0 : boolean;
  signal type_cast_2186_inst_req_1 : boolean;
  signal type_cast_2184_inst_req_1 : boolean;
  signal ptr_deref_2283_load_0_req_1 : boolean;
  signal ptr_deref_2283_load_0_ack_1 : boolean;
  signal phi_stmt_2174_req_0 : boolean;
  signal type_cast_2177_inst_ack_1 : boolean;
  signal phi_stmt_2181_ack_0 : boolean;
  signal type_cast_2287_inst_req_0 : boolean;
  signal type_cast_2287_inst_ack_0 : boolean;
  signal type_cast_2287_inst_req_1 : boolean;
  signal type_cast_2287_inst_ack_1 : boolean;
  signal array_obj_ref_2299_index_offset_req_0 : boolean;
  signal array_obj_ref_2299_index_offset_ack_0 : boolean;
  signal array_obj_ref_2299_index_offset_req_1 : boolean;
  signal array_obj_ref_2299_index_offset_ack_1 : boolean;
  signal addr_of_2300_final_reg_req_0 : boolean;
  signal addr_of_2300_final_reg_ack_0 : boolean;
  signal addr_of_2300_final_reg_req_1 : boolean;
  signal addr_of_2300_final_reg_ack_1 : boolean;
  signal ptr_deref_2303_store_0_req_0 : boolean;
  signal ptr_deref_2303_store_0_ack_0 : boolean;
  signal ptr_deref_2303_store_0_req_1 : boolean;
  signal ptr_deref_2303_store_0_ack_1 : boolean;
  signal type_cast_2308_inst_req_0 : boolean;
  signal type_cast_2308_inst_ack_0 : boolean;
  signal type_cast_2308_inst_req_1 : boolean;
  signal type_cast_2308_inst_ack_1 : boolean;
  signal if_stmt_2321_branch_req_0 : boolean;
  signal if_stmt_2321_branch_ack_1 : boolean;
  signal if_stmt_2321_branch_ack_0 : boolean;
  signal type_cast_2344_inst_req_0 : boolean;
  signal type_cast_2344_inst_ack_0 : boolean;
  signal type_cast_2344_inst_req_1 : boolean;
  signal type_cast_2344_inst_ack_1 : boolean;
  signal type_cast_2353_inst_req_0 : boolean;
  signal type_cast_2353_inst_ack_0 : boolean;
  signal type_cast_2353_inst_req_1 : boolean;
  signal type_cast_2353_inst_ack_1 : boolean;
  signal if_stmt_2372_branch_req_0 : boolean;
  signal if_stmt_2372_branch_ack_1 : boolean;
  signal if_stmt_2372_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2380_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2380_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2380_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2380_inst_ack_1 : boolean;
  signal phi_stmt_2174_req_1 : boolean;
  signal type_cast_2186_inst_req_0 : boolean;
  signal type_cast_2186_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5963_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5963_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5963_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5963_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5963: Block -- control-path 
    signal convTransposeC_CP_5963_elements: BooleanArray(79 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5963_elements(0) <= convTransposeC_CP_5963_start;
    convTransposeC_CP_5963_symbol <= convTransposeC_CP_5963_elements(57);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2018/assign_stmt_2021/$entry
      -- CP-element group 0: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2018/$entry
      -- CP-element group 0: 	 branch_block_stmt_2018/branch_block_stmt_2018__entry__
      -- CP-element group 0: 	 branch_block_stmt_2018/assign_stmt_2021__entry__
      -- 
    rr_6011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(0), ack => RPIPE_Block2_start_2020_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Update/$entry
      -- 
    ra_6012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2020_inst_ack_0, ack => convTransposeC_CP_5963_elements(1)); -- 
    cr_6016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(1), ack => RPIPE_Block2_start_2020_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (259) 
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2021/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2021/RPIPE_Block2_start_2020_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2021__exit__
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171__entry__
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Update/cr
      -- 
    ca_6017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2020_inst_ack_1, ack => convTransposeC_CP_5963_elements(2)); -- 
    cr_6064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2033_load_0_req_1); -- 
    rr_6053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2033_load_0_req_0); -- 
    rr_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2051_load_0_req_0); -- 
    cr_6114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2051_load_0_req_1); -- 
    rr_6153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2063_load_0_req_0); -- 
    cr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2063_load_0_req_1); -- 
    rr_6203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2073_load_0_req_0); -- 
    cr_6214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2073_load_0_req_1); -- 
    rr_6253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2085_load_0_req_0); -- 
    cr_6264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2085_load_0_req_1); -- 
    rr_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => LOAD_padding_2088_load_0_req_0); -- 
    cr_6297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => LOAD_padding_2088_load_0_req_1); -- 
    rr_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2098_load_0_req_0); -- 
    cr_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2098_load_0_req_1); -- 
    rr_6386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2110_load_0_req_0); -- 
    cr_6397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2110_load_0_req_1); -- 
    rr_6436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2122_load_0_req_0); -- 
    cr_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2122_load_0_req_1); -- 
    rr_6486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2134_load_0_req_0); -- 
    cr_6497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => ptr_deref_2134_load_0_req_1); -- 
    cr_6516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => type_cast_2138_inst_req_1); -- 
    cr_6530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(2), ack => type_cast_2142_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_sample_completed_
      -- 
    ra_6054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2033_load_0_ack_0, ack => convTransposeC_CP_5963_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/ptr_deref_2033_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/ptr_deref_2033_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/ptr_deref_2033_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2033_Update/ptr_deref_2033_Merge/merge_ack
      -- 
    ca_6065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2033_load_0_ack_1, ack => convTransposeC_CP_5963_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Sample/word_access_start/$exit
      -- 
    ra_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2051_load_0_ack_0, ack => convTransposeC_CP_5963_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/ptr_deref_2051_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/ptr_deref_2051_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/ptr_deref_2051_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2051_Update/ptr_deref_2051_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Sample/rr
      -- 
    ca_6115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2051_load_0_ack_1, ack => convTransposeC_CP_5963_elements(6)); -- 
    rr_6511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(6), ack => type_cast_2138_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Sample/word_access_start/word_0/ra
      -- 
    ra_6154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2063_load_0_ack_0, ack => convTransposeC_CP_5963_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	25 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/ptr_deref_2063_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/ptr_deref_2063_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/ptr_deref_2063_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2063_Update/ptr_deref_2063_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Sample/rr
      -- 
    ca_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2063_load_0_ack_1, ack => convTransposeC_CP_5963_elements(8)); -- 
    rr_6525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(8), ack => type_cast_2142_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Sample/word_access_start/word_0/ra
      -- 
    ra_6204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_load_0_ack_0, ack => convTransposeC_CP_5963_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	27 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/ptr_deref_2073_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/ptr_deref_2073_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/ptr_deref_2073_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2073_Update/ptr_deref_2073_Merge/merge_ack
      -- 
    ca_6215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2073_load_0_ack_1, ack => convTransposeC_CP_5963_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Sample/word_access_start/word_0/ra
      -- 
    ra_6254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2085_load_0_ack_0, ack => convTransposeC_CP_5963_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	27 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/ptr_deref_2085_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/ptr_deref_2085_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/ptr_deref_2085_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2085_Update/ptr_deref_2085_Merge/merge_ack
      -- 
    ca_6265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2085_load_0_ack_1, ack => convTransposeC_CP_5963_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Sample/word_access_start/word_0/ra
      -- 
    ra_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2088_load_0_ack_0, ack => convTransposeC_CP_5963_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/LOAD_padding_2088_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/LOAD_padding_2088_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/LOAD_padding_2088_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/LOAD_padding_2088_Update/LOAD_padding_2088_Merge/merge_ack
      -- 
    ca_6298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2088_load_0_ack_1, ack => convTransposeC_CP_5963_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Sample/word_access_start/word_0/ra
      -- 
    ra_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2098_load_0_ack_0, ack => convTransposeC_CP_5963_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	27 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/ptr_deref_2098_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/ptr_deref_2098_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/ptr_deref_2098_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2098_Update/ptr_deref_2098_Merge/merge_ack
      -- 
    ca_6348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2098_load_0_ack_1, ack => convTransposeC_CP_5963_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Sample/word_access_start/word_0/ra
      -- 
    ra_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_load_0_ack_0, ack => convTransposeC_CP_5963_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	27 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/ptr_deref_2110_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/ptr_deref_2110_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/ptr_deref_2110_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2110_Update/ptr_deref_2110_Merge/merge_ack
      -- 
    ca_6398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_load_0_ack_1, ack => convTransposeC_CP_5963_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Sample/word_access_start/word_0/ra
      -- 
    ra_6437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2122_load_0_ack_0, ack => convTransposeC_CP_5963_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	27 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/ptr_deref_2122_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/ptr_deref_2122_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/ptr_deref_2122_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2122_Update/ptr_deref_2122_Merge/merge_ack
      -- 
    ca_6448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2122_load_0_ack_1, ack => convTransposeC_CP_5963_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Sample/word_access_start/word_0/ra
      -- 
    ra_6487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2134_load_0_ack_0, ack => convTransposeC_CP_5963_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/ptr_deref_2134_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/ptr_deref_2134_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/ptr_deref_2134_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/ptr_deref_2134_Update/ptr_deref_2134_Merge/merge_ack
      -- 
    ca_6498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2134_load_0_ack_1, ack => convTransposeC_CP_5963_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Sample/ra
      -- 
    ra_6512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2138_inst_ack_0, ack => convTransposeC_CP_5963_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2138_Update/ca
      -- 
    ca_6517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2138_inst_ack_1, ack => convTransposeC_CP_5963_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	8 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Sample/ra
      -- 
    ra_6526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2142_inst_ack_0, ack => convTransposeC_CP_5963_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/type_cast_2142_Update/ca
      -- 
    ca_6531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2142_inst_ack_1, ack => convTransposeC_CP_5963_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  place  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	20 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	12 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	16 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	58 
    -- CP-element group 27: 	59 
    -- CP-element group 27: 	60 
    -- CP-element group 27:  members (14) 
      -- CP-element group 27: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171/$exit
      -- CP-element group 27: 	 branch_block_stmt_2018/assign_stmt_2030_to_assign_stmt_2171__exit__
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Update/cr
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Update/$entry
      -- 
    cr_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(27), ack => type_cast_2186_inst_req_1); -- 
    rr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(27), ack => type_cast_2186_inst_req_0); -- 
    convTransposeC_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(20) & convTransposeC_CP_5963_elements(22) & convTransposeC_CP_5963_elements(26) & convTransposeC_CP_5963_elements(24) & convTransposeC_CP_5963_elements(10) & convTransposeC_CP_5963_elements(12) & convTransposeC_CP_5963_elements(14) & convTransposeC_CP_5963_elements(16) & convTransposeC_CP_5963_elements(18) & convTransposeC_CP_5963_elements(4);
      gj_convTransposeC_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	79 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Sample/ra
      -- 
    ra_6546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_0, ack => convTransposeC_CP_5963_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	79 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (16) 
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Sample/req
      -- 
    ca_6551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_1, ack => convTransposeC_CP_5963_elements(29)); -- 
    req_6576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(29), ack => array_obj_ref_2278_index_offset_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	47 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_sample_complete
      -- CP-element group 30: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Sample/ack
      -- 
    ack_6577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2278_index_offset_ack_0, ack => convTransposeC_CP_5963_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	79 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (11) 
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_offset_calculated
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_request/$entry
      -- CP-element group 31: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_request/req
      -- 
    ack_6582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2278_index_offset_ack_1, ack => convTransposeC_CP_5963_elements(31)); -- 
    req_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(31), ack => addr_of_2279_final_reg_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_request/$exit
      -- CP-element group 32: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_request/ack
      -- 
    ack_6592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2279_final_reg_ack_0, ack => convTransposeC_CP_5963_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	79 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (24) 
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_complete/ack
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_word_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_address_resized
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_addr_resize/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_addr_resize/$exit
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_addr_resize/base_resize_req
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_addr_resize/base_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_word_addrgen/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_word_addrgen/$exit
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_word_addrgen/root_register_req
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_word_addrgen/root_register_ack
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/word_0/rr
      -- 
    ack_6597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2279_final_reg_ack_1, ack => convTransposeC_CP_5963_elements(33)); -- 
    rr_6630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(33), ack => ptr_deref_2283_load_0_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Sample/word_access_start/word_0/ra
      -- 
    ra_6631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_load_0_ack_0, ack => convTransposeC_CP_5963_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	79 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	42 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/ptr_deref_2283_Merge/$entry
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/ptr_deref_2283_Merge/$exit
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/ptr_deref_2283_Merge/merge_req
      -- CP-element group 35: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/ptr_deref_2283_Merge/merge_ack
      -- 
    ca_6642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2283_load_0_ack_1, ack => convTransposeC_CP_5963_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	79 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Sample/ra
      -- 
    ra_6656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_0, ack => convTransposeC_CP_5963_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	79 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Sample/req
      -- 
    ca_6661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2287_inst_ack_1, ack => convTransposeC_CP_5963_elements(37)); -- 
    req_6686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(37), ack => array_obj_ref_2299_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Sample/ack
      -- 
    ack_6687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2299_index_offset_ack_0, ack => convTransposeC_CP_5963_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	79 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_request/req
      -- 
    ack_6692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2299_index_offset_ack_1, ack => convTransposeC_CP_5963_elements(39)); -- 
    req_6701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(39), ack => addr_of_2300_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_request/ack
      -- 
    ack_6702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2300_final_reg_ack_0, ack => convTransposeC_CP_5963_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	79 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (19) 
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_word_addrgen/root_register_ack
      -- 
    ack_6707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2300_final_reg_ack_1, ack => convTransposeC_CP_5963_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	35 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/ptr_deref_2303_Split/$entry
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/ptr_deref_2303_Split/$exit
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/ptr_deref_2303_Split/split_req
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/ptr_deref_2303_Split/split_ack
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/word_0/rr
      -- 
    rr_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(42), ack => ptr_deref_2303_store_0_req_0); -- 
    convTransposeC_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(35) & convTransposeC_CP_5963_elements(41);
      gj_convTransposeC_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Sample/word_access_start/word_0/ra
      -- 
    ra_6746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2303_store_0_ack_0, ack => convTransposeC_CP_5963_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	79 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/word_0/ca
      -- 
    ca_6757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2303_store_0_ack_1, ack => convTransposeC_CP_5963_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	79 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Sample/ra
      -- 
    ra_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_0, ack => convTransposeC_CP_5963_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	79 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Update/ca
      -- 
    ca_6771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_1, ack => convTransposeC_CP_5963_elements(46)); -- 
    -- CP-element group 47:  branch  join  transition  place  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	30 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (10) 
      -- CP-element group 47: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320__exit__
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321__entry__
      -- CP-element group 47: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/$exit
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_2018/R_cmp_2322_place
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2018/if_stmt_2321_else_link/$entry
      -- 
    branch_req_6779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(47), ack => if_stmt_2321_branch_req_0); -- 
    convTransposeC_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(30) & convTransposeC_CP_5963_elements(44) & convTransposeC_CP_5963_elements(46) & convTransposeC_CP_5963_elements(38);
      gj_convTransposeC_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48: 	75 
    -- CP-element group 48:  members (24) 
      -- CP-element group 48: 	 branch_block_stmt_2018/merge_stmt_2327_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_2018/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_2018/merge_stmt_2327_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/merge_stmt_2327_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_2018/merge_stmt_2327_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_2018/merge_stmt_2327__exit__
      -- CP-element group 48: 	 branch_block_stmt_2018/assign_stmt_2333__entry__
      -- CP-element group 48: 	 branch_block_stmt_2018/assign_stmt_2333__exit__
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/cr
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/if_stmt_2321_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_2018/if_stmt_2321_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_2018/whilex_xbody_ifx_xthen
      -- CP-element group 48: 	 branch_block_stmt_2018/assign_stmt_2333/$entry
      -- CP-element group 48: 	 branch_block_stmt_2018/assign_stmt_2333/$exit
      -- 
    if_choice_transition_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2321_branch_ack_1, ack => convTransposeC_CP_5963_elements(48)); -- 
    cr_6973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(48), ack => type_cast_2243_inst_req_1); -- 
    rr_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(48), ack => type_cast_2243_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	53 
    -- CP-element group 49:  members (21) 
      -- CP-element group 49: 	 branch_block_stmt_2018/merge_stmt_2335_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_2018/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/merge_stmt_2335__exit__
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371__entry__
      -- CP-element group 49: 	 branch_block_stmt_2018/merge_stmt_2335_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_2018/merge_stmt_2335_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_2018/merge_stmt_2335_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_2018/if_stmt_2321_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_2018/if_stmt_2321_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_2018/whilex_xbody_ifx_xelse
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_update_start_
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_update_start_
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Update/cr
      -- 
    else_choice_transition_6788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2321_branch_ack_0, ack => convTransposeC_CP_5963_elements(49)); -- 
    rr_6804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(49), ack => type_cast_2344_inst_req_0); -- 
    cr_6809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(49), ack => type_cast_2344_inst_req_1); -- 
    cr_6823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(49), ack => type_cast_2353_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Sample/ra
      -- 
    ra_6805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_0, ack => convTransposeC_CP_5963_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2344_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Sample/rr
      -- 
    ca_6810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2344_inst_ack_1, ack => convTransposeC_CP_5963_elements(51)); -- 
    rr_6818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(51), ack => type_cast_2353_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Sample/ra
      -- 
    ra_6819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_0, ack => convTransposeC_CP_5963_elements(52)); -- 
    -- CP-element group 53:  branch  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	49 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (13) 
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372__entry__
      -- CP-element group 53: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371__exit__
      -- CP-element group 53: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/$exit
      -- CP-element group 53: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2018/assign_stmt_2341_to_assign_stmt_2371/type_cast_2353_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_2018/R_cmp97_2373_place
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2018/if_stmt_2372_else_link/$entry
      -- 
    ca_6824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2353_inst_ack_1, ack => convTransposeC_CP_5963_elements(53)); -- 
    branch_req_6832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(53), ack => if_stmt_2372_branch_req_0); -- 
    -- CP-element group 54:  merge  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (15) 
      -- CP-element group 54: 	 branch_block_stmt_2018/merge_stmt_2378__exit__
      -- CP-element group 54: 	 branch_block_stmt_2018/merge_stmt_2378_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_2018/assign_stmt_2382__entry__
      -- CP-element group 54: 	 branch_block_stmt_2018/merge_stmt_2378_PhiAck/dummy
      -- CP-element group 54: 	 branch_block_stmt_2018/merge_stmt_2378_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_2018/merge_stmt_2378_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_2018/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_2018/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2018/if_stmt_2372_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_2018/if_stmt_2372_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_2018/ifx_xelse_whilex_xend
      -- CP-element group 54: 	 branch_block_stmt_2018/assign_stmt_2382/$entry
      -- CP-element group 54: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Sample/req
      -- 
    if_choice_transition_6837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2372_branch_ack_1, ack => convTransposeC_CP_5963_elements(54)); -- 
    req_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(54), ack => WPIPE_Block2_done_2380_inst_req_0); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	63 
    -- CP-element group 55: 	64 
    -- CP-element group 55: 	66 
    -- CP-element group 55: 	67 
    -- CP-element group 55:  members (20) 
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2018/if_stmt_2372_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2018/if_stmt_2372_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter
      -- 
    else_choice_transition_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2372_branch_ack_0, ack => convTransposeC_CP_5963_elements(55)); -- 
    rr_6913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(55), ack => type_cast_2177_inst_req_0); -- 
    rr_6936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(55), ack => type_cast_2184_inst_req_0); -- 
    cr_6918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(55), ack => type_cast_2177_inst_req_1); -- 
    cr_6941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(55), ack => type_cast_2184_inst_req_1); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Update/req
      -- 
    ack_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2380_inst_ack_0, ack => convTransposeC_CP_5963_elements(56)); -- 
    req_6859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(56), ack => WPIPE_Block2_done_2380_inst_req_1); -- 
    -- CP-element group 57:  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (16) 
      -- CP-element group 57: 	 branch_block_stmt_2018/merge_stmt_2384_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2018/assign_stmt_2382__exit__
      -- CP-element group 57: 	 branch_block_stmt_2018/return__
      -- CP-element group 57: 	 branch_block_stmt_2018/merge_stmt_2384__exit__
      -- CP-element group 57: 	 $exit
      -- CP-element group 57: 	 branch_block_stmt_2018/$exit
      -- CP-element group 57: 	 branch_block_stmt_2018/branch_block_stmt_2018__exit__
      -- CP-element group 57: 	 branch_block_stmt_2018/merge_stmt_2384_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_2018/merge_stmt_2384_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2018/merge_stmt_2384_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2018/return___PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2018/return___PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_2018/assign_stmt_2382/$exit
      -- CP-element group 57: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2018/assign_stmt_2382/WPIPE_Block2_done_2380_Update/ack
      -- 
    ack_6860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2380_inst_ack_1, ack => convTransposeC_CP_5963_elements(57)); -- 
    -- CP-element group 58:  transition  output  delay-element  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	27 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	62 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/$exit
      -- CP-element group 58: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/$exit
      -- CP-element group 58: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2180_konst_delay_trans
      -- CP-element group 58: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_req
      -- 
    phi_stmt_2174_req_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2174_req_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(58), ack => phi_stmt_2174_req_1); -- 
    -- Element group convTransposeC_CP_5963_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => convTransposeC_CP_5963_elements(27), ack => convTransposeC_CP_5963_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	27 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Sample/ra
      -- 
    ra_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_0, ack => convTransposeC_CP_5963_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Update/ca
      -- CP-element group 60: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/Update/$exit
      -- 
    ca_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_1, ack => convTransposeC_CP_5963_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_req
      -- CP-element group 61: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/$exit
      -- CP-element group 61: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$exit
      -- CP-element group 61: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/$exit
      -- CP-element group 61: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2186/SplitProtocol/$exit
      -- 
    phi_stmt_2181_req_6894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2181_req_6894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(61), ack => phi_stmt_2181_req_1); -- 
    convTransposeC_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(59) & convTransposeC_CP_5963_elements(60);
      gj_convTransposeC_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	70 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_2018/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(58) & convTransposeC_CP_5963_elements(61);
      gj_convTransposeC_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	55 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Sample/$exit
      -- 
    ra_6914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2177_inst_ack_0, ack => convTransposeC_CP_5963_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	55 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/Update/ca
      -- 
    ca_6919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2177_inst_ack_1, ack => convTransposeC_CP_5963_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	69 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/$exit
      -- CP-element group 65: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/$exit
      -- CP-element group 65: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_sources/type_cast_2177/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2174/phi_stmt_2174_req
      -- 
    phi_stmt_2174_req_6920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2174_req_6920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(65), ack => phi_stmt_2174_req_0); -- 
    convTransposeC_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(63) & convTransposeC_CP_5963_elements(64);
      gj_convTransposeC_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	55 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Sample/ra
      -- 
    ra_6937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_0, ack => convTransposeC_CP_5963_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	55 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/Update/ca
      -- 
    ca_6942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_1, ack => convTransposeC_CP_5963_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/$exit
      -- CP-element group 68: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/type_cast_2184/SplitProtocol/$exit
      -- CP-element group 68: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/$exit
      -- CP-element group 68: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2181/phi_stmt_2181_req
      -- 
    phi_stmt_2181_req_6943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2181_req_6943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(68), ack => phi_stmt_2181_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(66) & convTransposeC_CP_5963_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	65 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2018/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(65) & convTransposeC_CP_5963_elements(68);
      gj_convTransposeC_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  merge  fork  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	62 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2018/merge_stmt_2173_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2018/merge_stmt_2173_PhiReqMerge
      -- 
    convTransposeC_CP_5963_elements(70) <= OrReduce(convTransposeC_CP_5963_elements(62) & convTransposeC_CP_5963_elements(69));
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2018/merge_stmt_2173_PhiAck/phi_stmt_2174_ack
      -- 
    phi_stmt_2174_ack_6948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2174_ack_0, ack => convTransposeC_CP_5963_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2018/merge_stmt_2173_PhiAck/phi_stmt_2181_ack
      -- 
    phi_stmt_2181_ack_6949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2181_ack_0, ack => convTransposeC_CP_5963_elements(72)); -- 
    -- CP-element group 73:  join  transition  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (10) 
      -- CP-element group 73: 	 branch_block_stmt_2018/merge_stmt_2173_PhiAck/$exit
      -- CP-element group 73: 	 branch_block_stmt_2018/merge_stmt_2173__exit__
      -- CP-element group 73: 	 branch_block_stmt_2018/assign_stmt_2192_to_assign_stmt_2237__entry__
      -- CP-element group 73: 	 branch_block_stmt_2018/assign_stmt_2192_to_assign_stmt_2237__exit__
      -- CP-element group 73: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 73: 	 branch_block_stmt_2018/assign_stmt_2192_to_assign_stmt_2237/$entry
      -- CP-element group 73: 	 branch_block_stmt_2018/assign_stmt_2192_to_assign_stmt_2237/$exit
      -- CP-element group 73: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/$entry
      -- CP-element group 73: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- 
    convTransposeC_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(71) & convTransposeC_CP_5963_elements(72);
      gj_convTransposeC_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	48 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Sample/$exit
      -- 
    ra_6969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_0, ack => convTransposeC_CP_5963_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	48 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/Update/$exit
      -- 
    ca_6974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2243_inst_ack_1, ack => convTransposeC_CP_5963_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2243/$exit
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 76: 	 branch_block_stmt_2018/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2240_req_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(76), ack => phi_stmt_2240_req_0); -- 
    convTransposeC_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5963_elements(74) & convTransposeC_CP_5963_elements(75);
      gj_convTransposeC_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5963_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_req
      -- CP-element group 77: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/type_cast_2246_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/phi_stmt_2240_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2240/$exit
      -- CP-element group 77: 	 branch_block_stmt_2018/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2240_req_6986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2240_req_6986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(77), ack => phi_stmt_2240_req_1); -- 
    -- Element group convTransposeC_CP_5963_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeC_CP_5963_elements(73), ack => convTransposeC_CP_5963_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  merge  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2018/merge_stmt_2239_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2018/merge_stmt_2239_PhiReqMerge
      -- 
    convTransposeC_CP_5963_elements(78) <= OrReduce(convTransposeC_CP_5963_elements(76) & convTransposeC_CP_5963_elements(77));
    -- CP-element group 79:  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	28 
    -- CP-element group 79: 	29 
    -- CP-element group 79: 	31 
    -- CP-element group 79: 	33 
    -- CP-element group 79: 	35 
    -- CP-element group 79: 	36 
    -- CP-element group 79: 	37 
    -- CP-element group 79: 	41 
    -- CP-element group 79: 	44 
    -- CP-element group 79: 	45 
    -- CP-element group 79: 	46 
    -- CP-element group 79: 	39 
    -- CP-element group 79:  members (45) 
      -- CP-element group 79: 	 branch_block_stmt_2018/merge_stmt_2239_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_2018/merge_stmt_2239_PhiAck/phi_stmt_2240_ack
      -- CP-element group 79: 	 branch_block_stmt_2018/merge_stmt_2239__exit__
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320__entry__
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2266_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_update_start
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2278_final_index_sum_regn_Update/req
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2279_complete/req
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/word_0/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2283_Update/word_access_complete/word_0/cr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2287_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_update_start
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/array_obj_ref_2299_final_index_sum_regn_Update/req
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/addr_of_2300_complete/req
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/word_0/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/ptr_deref_2303_Update/word_access_complete/word_0/cr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2018/assign_stmt_2253_to_assign_stmt_2320/type_cast_2308_Update/cr
      -- 
    phi_stmt_2240_ack_6991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2240_ack_0, ack => convTransposeC_CP_5963_elements(79)); -- 
    rr_6545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2266_inst_req_0); -- 
    cr_6550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2266_inst_req_1); -- 
    req_6581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => array_obj_ref_2278_index_offset_req_1); -- 
    req_6596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => addr_of_2279_final_reg_req_1); -- 
    cr_6641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => ptr_deref_2283_load_0_req_1); -- 
    rr_6655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2287_inst_req_0); -- 
    cr_6660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2287_inst_req_1); -- 
    req_6691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => array_obj_ref_2299_index_offset_req_1); -- 
    req_6706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => addr_of_2300_final_reg_req_1); -- 
    cr_6756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => ptr_deref_2303_store_0_req_1); -- 
    rr_6765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2308_inst_req_0); -- 
    cr_6770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5963_elements(79), ack => type_cast_2308_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_2088_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2088_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr111_2277_resized : std_logic_vector(13 downto 0);
    signal R_shr111_2277_scaled : std_logic_vector(13 downto 0);
    signal R_shr68113_2298_resized : std_logic_vector(13 downto 0);
    signal R_shr68113_2298_scaled : std_logic_vector(13 downto 0);
    signal add21_2258 : std_logic_vector(15 downto 0);
    signal add61_2263 : std_logic_vector(15 downto 0);
    signal add74_2315 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2278_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2278_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2278_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2278_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2278_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2278_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2299_root_address : std_logic_vector(13 downto 0);
    signal arrayidx70_2301 : std_logic_vector(31 downto 0);
    signal arrayidx_2280 : std_logic_vector(31 downto 0);
    signal call_2021 : std_logic_vector(15 downto 0);
    signal cmp88_2350 : std_logic_vector(0 downto 0);
    signal cmp97_2371 : std_logic_vector(0 downto 0);
    signal cmp_2320 : std_logic_vector(0 downto 0);
    signal conv64_2267 : std_logic_vector(63 downto 0);
    signal conv67_2288 : std_logic_vector(63 downto 0);
    signal conv73_2309 : std_logic_vector(31 downto 0);
    signal conv76_2139 : std_logic_vector(31 downto 0);
    signal conv84_2345 : std_logic_vector(31 downto 0);
    signal conv86_2143 : std_logic_vector(31 downto 0);
    signal div87_2149 : std_logic_vector(31 downto 0);
    signal div_2040 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2131 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2030 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2048 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2060 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2070 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2082 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2095 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2107 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2119 : std_logic_vector(31 downto 0);
    signal inc92_2354 : std_logic_vector(15 downto 0);
    signal inc92x_xinput_dim0x_x2_2359 : std_logic_vector(15 downto 0);
    signal inc_2341 : std_logic_vector(15 downto 0);
    signal indvar_2240 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2333 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2181 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2174 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2366 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2253 : std_logic_vector(15 downto 0);
    signal ptr_deref_2033_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2033_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2033_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2033_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2033_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2051_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2051_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2051_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2051_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2051_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2063_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2063_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2063_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2063_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2063_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2073_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2073_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2073_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2073_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2073_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2085_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2085_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2085_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2085_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2085_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2098_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2098_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2098_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2098_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2098_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2110_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2110_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2110_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2110_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2110_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2122_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2122_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2122_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2122_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2122_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2134_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2134_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2134_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2134_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2134_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2283_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2283_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2283_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2283_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2283_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2303_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2303_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2303_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2303_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2303_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2303_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr111_2273 : std_logic_vector(63 downto 0);
    signal shr68113_2294 : std_logic_vector(63 downto 0);
    signal tmp10_2222 : std_logic_vector(15 downto 0);
    signal tmp11_2227 : std_logic_vector(15 downto 0);
    signal tmp127_2192 : std_logic_vector(15 downto 0);
    signal tmp128_2197 : std_logic_vector(15 downto 0);
    signal tmp129_2202 : std_logic_vector(15 downto 0);
    signal tmp12_2052 : std_logic_vector(15 downto 0);
    signal tmp13_2232 : std_logic_vector(15 downto 0);
    signal tmp14_2237 : std_logic_vector(15 downto 0);
    signal tmp16_2064 : std_logic_vector(15 downto 0);
    signal tmp25_2074 : std_logic_vector(15 downto 0);
    signal tmp28_2086 : std_logic_vector(15 downto 0);
    signal tmp31_2089 : std_logic_vector(15 downto 0);
    signal tmp37_2099 : std_logic_vector(15 downto 0);
    signal tmp3_2155 : std_logic_vector(15 downto 0);
    signal tmp40_2111 : std_logic_vector(15 downto 0);
    signal tmp4_2160 : std_logic_vector(15 downto 0);
    signal tmp50_2123 : std_logic_vector(15 downto 0);
    signal tmp54_2135 : std_logic_vector(15 downto 0);
    signal tmp5_2207 : std_logic_vector(15 downto 0);
    signal tmp65_2284 : std_logic_vector(63 downto 0);
    signal tmp6_2212 : std_logic_vector(15 downto 0);
    signal tmp7_2166 : std_logic_vector(15 downto 0);
    signal tmp8_2171 : std_logic_vector(15 downto 0);
    signal tmp9_2217 : std_logic_vector(15 downto 0);
    signal tmp_2034 : std_logic_vector(15 downto 0);
    signal type_cast_2038_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2147_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2153_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2164_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2177_wire : std_logic_vector(15 downto 0);
    signal type_cast_2180_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2184_wire : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire : std_logic_vector(15 downto 0);
    signal type_cast_2243_wire : std_logic_vector(15 downto 0);
    signal type_cast_2246_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2271_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2292_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2313_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2331_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2339_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2363_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_2088_word_address_0 <= "0";
    array_obj_ref_2278_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2278_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2278_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2278_resized_base_address <= "00000000000000";
    array_obj_ref_2299_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2299_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2299_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2299_resized_base_address <= "00000000000000";
    iNsTr_10_2131 <= "00000000000000000000000000000100";
    iNsTr_2_2030 <= "00000000000000000000000000000011";
    iNsTr_3_2048 <= "00000000000000000000000000000101";
    iNsTr_4_2060 <= "00000000000000000000000000000100";
    iNsTr_5_2070 <= "00000000000000000000000000000000";
    iNsTr_6_2082 <= "00000000000000000000000000000100";
    iNsTr_7_2095 <= "00000000000000000000000000000001";
    iNsTr_8_2107 <= "00000000000000000000000000000101";
    iNsTr_9_2119 <= "00000000000000000000000000000101";
    ptr_deref_2033_word_offset_0 <= "0000000";
    ptr_deref_2051_word_offset_0 <= "0000000";
    ptr_deref_2063_word_offset_0 <= "0000000";
    ptr_deref_2073_word_offset_0 <= "0";
    ptr_deref_2085_word_offset_0 <= "0000000";
    ptr_deref_2098_word_offset_0 <= "0";
    ptr_deref_2110_word_offset_0 <= "0000000";
    ptr_deref_2122_word_offset_0 <= "0000000";
    ptr_deref_2134_word_offset_0 <= "0000000";
    ptr_deref_2283_word_offset_0 <= "00000000000000";
    ptr_deref_2303_word_offset_0 <= "00000000000000";
    type_cast_2038_wire_constant <= "0000000000000001";
    type_cast_2147_wire_constant <= "00000000000000000000000000000001";
    type_cast_2153_wire_constant <= "1111111111111111";
    type_cast_2164_wire_constant <= "1111111111111111";
    type_cast_2180_wire_constant <= "0000000000000000";
    type_cast_2246_wire_constant <= "0000000000000000";
    type_cast_2251_wire_constant <= "0000000000000100";
    type_cast_2271_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2292_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2313_wire_constant <= "00000000000000000000000000000100";
    type_cast_2331_wire_constant <= "0000000000000001";
    type_cast_2339_wire_constant <= "0000000000000001";
    type_cast_2363_wire_constant <= "0000000000000000";
    phi_stmt_2174: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2177_wire & type_cast_2180_wire_constant;
      req <= phi_stmt_2174_req_0 & phi_stmt_2174_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2174",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2174_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2174,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2174
    phi_stmt_2181: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2184_wire & type_cast_2186_wire;
      req <= phi_stmt_2181_req_0 & phi_stmt_2181_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2181",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2181_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2181,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2181
    phi_stmt_2240: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2243_wire & type_cast_2246_wire_constant;
      req <= phi_stmt_2240_req_0 & phi_stmt_2240_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2240",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2240_ack_0,
          idata => idata,
          odata => indvar_2240,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2240
    -- flow-through select operator MUX_2365_inst
    input_dim1x_x2_2366 <= type_cast_2363_wire_constant when (cmp88_2350(0) /=  '0') else inc_2341;
    addr_of_2279_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2279_final_reg_req_0;
      addr_of_2279_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2279_final_reg_req_1;
      addr_of_2279_final_reg_ack_1<= rack(0);
      addr_of_2279_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2279_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2278_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2300_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2300_final_reg_req_0;
      addr_of_2300_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2300_final_reg_req_1;
      addr_of_2300_final_reg_ack_1<= rack(0);
      addr_of_2300_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2300_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2299_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx70_2301,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2138_inst_req_0;
      type_cast_2138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2138_inst_req_1;
      type_cast_2138_inst_ack_1<= rack(0);
      type_cast_2138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_2052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2142_inst_req_0;
      type_cast_2142_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2142_inst_req_1;
      type_cast_2142_inst_ack_1<= rack(0);
      type_cast_2142_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2142_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2064,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2143,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2177_inst_req_0;
      type_cast_2177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2177_inst_req_1;
      type_cast_2177_inst_ack_1<= rack(0);
      type_cast_2177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2177_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2184_inst_req_0;
      type_cast_2184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2184_inst_req_1;
      type_cast_2184_inst_ack_1<= rack(0);
      type_cast_2184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc92x_xinput_dim0x_x2_2359,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2184_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2186_inst_req_0;
      type_cast_2186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2186_inst_req_1;
      type_cast_2186_inst_ack_1<= rack(0);
      type_cast_2186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2040,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2243_inst_req_0;
      type_cast_2243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2243_inst_req_1;
      type_cast_2243_inst_ack_1<= rack(0);
      type_cast_2243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2243_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2266_inst_req_0;
      type_cast_2266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2266_inst_req_1;
      type_cast_2266_inst_ack_1<= rack(0);
      type_cast_2266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_2258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_2267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2287_inst_req_0;
      type_cast_2287_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2287_inst_req_1;
      type_cast_2287_inst_ack_1<= rack(0);
      type_cast_2287_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2287_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add61_2263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_2288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2308_inst_req_0;
      type_cast_2308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2308_inst_req_1;
      type_cast_2308_inst_ack_1<= rack(0);
      type_cast_2308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2344_inst_req_0;
      type_cast_2344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2344_inst_req_1;
      type_cast_2344_inst_ack_1<= rack(0);
      type_cast_2344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2345,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2353_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2353_inst_req_0;
      type_cast_2353_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2353_inst_req_1;
      type_cast_2353_inst_ack_1<= rack(0);
      type_cast_2353_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2353_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp88_2350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc92_2354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2088_gather_scatter
    process(LOAD_padding_2088_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2088_data_0;
      ov(15 downto 0) := iv;
      tmp31_2089 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2278_index_1_rename
    process(R_shr111_2277_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr111_2277_resized;
      ov(13 downto 0) := iv;
      R_shr111_2277_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2278_index_1_resize
    process(shr111_2273) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr111_2273;
      ov := iv(13 downto 0);
      R_shr111_2277_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2278_root_address_inst
    process(array_obj_ref_2278_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2278_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2278_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2299_index_1_rename
    process(R_shr68113_2298_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr68113_2298_resized;
      ov(13 downto 0) := iv;
      R_shr68113_2298_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2299_index_1_resize
    process(shr68113_2294) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr68113_2294;
      ov := iv(13 downto 0);
      R_shr68113_2298_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2299_root_address_inst
    process(array_obj_ref_2299_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2299_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2299_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2033_addr_0
    process(ptr_deref_2033_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2033_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2033_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2033_base_resize
    process(iNsTr_2_2030) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2030;
      ov := iv(6 downto 0);
      ptr_deref_2033_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2033_gather_scatter
    process(ptr_deref_2033_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2033_data_0;
      ov(15 downto 0) := iv;
      tmp_2034 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2033_root_address_inst
    process(ptr_deref_2033_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2033_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2033_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2051_addr_0
    process(ptr_deref_2051_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2051_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2051_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2051_base_resize
    process(iNsTr_3_2048) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2048;
      ov := iv(6 downto 0);
      ptr_deref_2051_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2051_gather_scatter
    process(ptr_deref_2051_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2051_data_0;
      ov(15 downto 0) := iv;
      tmp12_2052 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2051_root_address_inst
    process(ptr_deref_2051_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2051_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2051_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2063_addr_0
    process(ptr_deref_2063_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2063_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2063_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2063_base_resize
    process(iNsTr_4_2060) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2060;
      ov := iv(6 downto 0);
      ptr_deref_2063_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2063_gather_scatter
    process(ptr_deref_2063_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2063_data_0;
      ov(15 downto 0) := iv;
      tmp16_2064 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2063_root_address_inst
    process(ptr_deref_2063_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2063_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2063_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_addr_0
    process(ptr_deref_2073_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2073_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_base_resize
    process(iNsTr_5_2070) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2070;
      ov := iv(0 downto 0);
      ptr_deref_2073_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_gather_scatter
    process(ptr_deref_2073_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_data_0;
      ov(15 downto 0) := iv;
      tmp25_2074 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2073_root_address_inst
    process(ptr_deref_2073_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2073_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2073_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2085_addr_0
    process(ptr_deref_2085_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2085_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2085_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2085_base_resize
    process(iNsTr_6_2082) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2082;
      ov := iv(6 downto 0);
      ptr_deref_2085_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2085_gather_scatter
    process(ptr_deref_2085_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2085_data_0;
      ov(15 downto 0) := iv;
      tmp28_2086 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2085_root_address_inst
    process(ptr_deref_2085_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2085_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2085_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2098_addr_0
    process(ptr_deref_2098_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2098_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2098_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2098_base_resize
    process(iNsTr_7_2095) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2095;
      ov := iv(0 downto 0);
      ptr_deref_2098_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2098_gather_scatter
    process(ptr_deref_2098_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2098_data_0;
      ov(15 downto 0) := iv;
      tmp37_2099 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2098_root_address_inst
    process(ptr_deref_2098_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2098_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2098_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2110_addr_0
    process(ptr_deref_2110_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2110_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2110_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2110_base_resize
    process(iNsTr_8_2107) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2107;
      ov := iv(6 downto 0);
      ptr_deref_2110_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2110_gather_scatter
    process(ptr_deref_2110_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2110_data_0;
      ov(15 downto 0) := iv;
      tmp40_2111 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2110_root_address_inst
    process(ptr_deref_2110_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2110_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2110_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2122_addr_0
    process(ptr_deref_2122_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2122_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2122_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2122_base_resize
    process(iNsTr_9_2119) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2119;
      ov := iv(6 downto 0);
      ptr_deref_2122_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2122_gather_scatter
    process(ptr_deref_2122_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2122_data_0;
      ov(15 downto 0) := iv;
      tmp50_2123 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2122_root_address_inst
    process(ptr_deref_2122_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2122_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2122_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_addr_0
    process(ptr_deref_2134_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2134_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2134_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_base_resize
    process(iNsTr_10_2131) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2131;
      ov := iv(6 downto 0);
      ptr_deref_2134_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_gather_scatter
    process(ptr_deref_2134_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2134_data_0;
      ov(15 downto 0) := iv;
      tmp54_2135 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2134_root_address_inst
    process(ptr_deref_2134_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2134_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2134_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2283_addr_0
    process(ptr_deref_2283_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2283_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2283_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2283_base_resize
    process(arrayidx_2280) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2280;
      ov := iv(13 downto 0);
      ptr_deref_2283_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2283_gather_scatter
    process(ptr_deref_2283_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2283_data_0;
      ov(63 downto 0) := iv;
      tmp65_2284 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2283_root_address_inst
    process(ptr_deref_2283_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2283_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2283_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2303_addr_0
    process(ptr_deref_2303_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2303_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2303_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2303_base_resize
    process(arrayidx70_2301) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx70_2301;
      ov := iv(13 downto 0);
      ptr_deref_2303_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2303_gather_scatter
    process(tmp65_2284) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp65_2284;
      ov(63 downto 0) := iv;
      ptr_deref_2303_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2303_root_address_inst
    process(ptr_deref_2303_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2303_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2303_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2320;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2321_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2321_branch_req_0,
          ack0 => if_stmt_2321_branch_ack_0,
          ack1 => if_stmt_2321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2372_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp97_2371;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2372_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2372_branch_req_0,
          ack0 => if_stmt_2372_branch_ack_0,
          ack1 => if_stmt_2372_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2154_inst
    process(tmp40_2111) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp40_2111, type_cast_2153_wire_constant, tmp_var);
      tmp3_2155 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2165_inst
    process(tmp28_2086) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp28_2086, type_cast_2164_wire_constant, tmp_var);
      tmp7_2166 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2196_inst
    process(input_dim1x_x1x_xph_2174, tmp127_2192) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2174, tmp127_2192, tmp_var);
      tmp128_2197 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2211_inst
    process(tmp4_2160, tmp5_2207) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_2160, tmp5_2207, tmp_var);
      tmp6_2212 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2221_inst
    process(tmp8_2171, tmp9_2217) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_2171, tmp9_2217, tmp_var);
      tmp10_2222 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2231_inst
    process(tmp6_2212, tmp11_2227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_2212, tmp11_2227, tmp_var);
      tmp13_2232 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2257_inst
    process(tmp129_2202, input_dim2x_x1_2253) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp129_2202, input_dim2x_x1_2253, tmp_var);
      add21_2258 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2262_inst
    process(tmp14_2237, input_dim2x_x1_2253) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2237, input_dim2x_x1_2253, tmp_var);
      add61_2263 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2332_inst
    process(indvar_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2240, type_cast_2331_wire_constant, tmp_var);
      indvarx_xnext_2333 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2340_inst
    process(input_dim1x_x1x_xph_2174) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2174, type_cast_2339_wire_constant, tmp_var);
      inc_2341 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2358_inst
    process(inc92_2354, input_dim0x_x2x_xph_2181) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc92_2354, input_dim0x_x2x_xph_2181, tmp_var);
      inc92x_xinput_dim0x_x2_2359 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2314_inst
    process(conv73_2309) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv73_2309, type_cast_2313_wire_constant, tmp_var);
      add74_2315 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2370_inst
    process(inc92x_xinput_dim0x_x2_2359, tmp_2034) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc92x_xinput_dim0x_x2_2359, tmp_2034, tmp_var);
      cmp97_2371 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2349_inst
    process(conv84_2345, div87_2149) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv84_2345, div87_2149, tmp_var);
      cmp88_2350 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2039_inst
    process(tmp_2034) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2034, type_cast_2038_wire_constant, tmp_var);
      div_2040 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2148_inst
    process(conv86_2143) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv86_2143, type_cast_2147_wire_constant, tmp_var);
      div87_2149 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2272_inst
    process(conv64_2267) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv64_2267, type_cast_2271_wire_constant, tmp_var);
      shr111_2273 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2293_inst
    process(conv67_2288) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv67_2288, type_cast_2292_wire_constant, tmp_var);
      shr68113_2294 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2191_inst
    process(tmp16_2064, input_dim0x_x2x_xph_2181) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2064, input_dim0x_x2x_xph_2181, tmp_var);
      tmp127_2192 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2201_inst
    process(tmp12_2052, tmp128_2197) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_2052, tmp128_2197, tmp_var);
      tmp129_2202 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2206_inst
    process(tmp37_2099, input_dim1x_x1x_xph_2174) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp37_2099, input_dim1x_x1x_xph_2174, tmp_var);
      tmp5_2207 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2216_inst
    process(tmp25_2074, input_dim0x_x2x_xph_2181) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_2074, input_dim0x_x2x_xph_2181, tmp_var);
      tmp9_2217 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2226_inst
    process(tmp54_2135, tmp10_2222) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_2135, tmp10_2222, tmp_var);
      tmp11_2227 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2236_inst
    process(tmp50_2123, tmp13_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp50_2123, tmp13_2232, tmp_var);
      tmp14_2237 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2252_inst
    process(indvar_2240) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2240, type_cast_2251_wire_constant, tmp_var);
      input_dim2x_x1_2253 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2159_inst
    process(tmp3_2155, tmp31_2089) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_2155, tmp31_2089, tmp_var);
      tmp4_2160 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2170_inst
    process(tmp7_2166, tmp31_2089) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_2166, tmp31_2089, tmp_var);
      tmp8_2171 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2319_inst
    process(add74_2315, conv76_2139) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add74_2315, conv76_2139, tmp_var);
      cmp_2320 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2278_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr111_2277_scaled;
      array_obj_ref_2278_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2278_index_offset_req_0;
      array_obj_ref_2278_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2278_index_offset_req_1;
      array_obj_ref_2278_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2299_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr68113_2298_scaled;
      array_obj_ref_2299_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2299_index_offset_req_0;
      array_obj_ref_2299_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2299_index_offset_req_1;
      array_obj_ref_2299_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : LOAD_padding_2088_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2088_load_0_req_0;
      LOAD_padding_2088_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2088_load_0_req_1;
      LOAD_padding_2088_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2088_word_address_0;
      LOAD_padding_2088_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2033_load_0 ptr_deref_2063_load_0 ptr_deref_2051_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2033_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2063_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2051_load_0_req_0;
      ptr_deref_2033_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2063_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2051_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2033_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2063_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2051_load_0_req_1;
      ptr_deref_2033_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2063_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2051_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2033_word_address_0 & ptr_deref_2063_word_address_0 & ptr_deref_2051_word_address_0;
      ptr_deref_2033_data_0 <= data_out(47 downto 32);
      ptr_deref_2063_data_0 <= data_out(31 downto 16);
      ptr_deref_2051_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2073_load_0 ptr_deref_2098_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2073_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2098_load_0_req_0;
      ptr_deref_2073_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2098_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2073_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2098_load_0_req_1;
      ptr_deref_2073_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2098_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2073_word_address_0 & ptr_deref_2098_word_address_0;
      ptr_deref_2073_data_0 <= data_out(31 downto 16);
      ptr_deref_2098_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2110_load_0 ptr_deref_2085_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2110_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2085_load_0_req_0;
      ptr_deref_2110_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2085_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2110_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2085_load_0_req_1;
      ptr_deref_2110_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2085_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2110_word_address_0 & ptr_deref_2085_word_address_0;
      ptr_deref_2110_data_0 <= data_out(31 downto 16);
      ptr_deref_2085_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2134_load_0 ptr_deref_2122_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2134_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2122_load_0_req_0;
      ptr_deref_2134_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2122_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2134_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2122_load_0_req_1;
      ptr_deref_2134_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2122_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2134_word_address_0 & ptr_deref_2122_word_address_0;
      ptr_deref_2134_data_0 <= data_out(31 downto 16);
      ptr_deref_2122_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2283_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2283_load_0_req_0;
      ptr_deref_2283_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2283_load_0_req_1;
      ptr_deref_2283_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2283_word_address_0;
      ptr_deref_2283_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2303_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2303_store_0_req_0;
      ptr_deref_2303_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2303_store_0_req_1;
      ptr_deref_2303_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2303_word_address_0;
      data_in <= ptr_deref_2303_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2020_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2020_inst_req_0;
      RPIPE_Block2_start_2020_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2020_inst_req_1;
      RPIPE_Block2_start_2020_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2021 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2380_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2380_inst_req_0;
      WPIPE_Block2_done_2380_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2380_inst_req_1;
      WPIPE_Block2_done_2380_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2021;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7032_start: Boolean;
  signal convTransposeD_CP_7032_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2611_inst_ack_0 : boolean;
  signal phi_stmt_2605_ack_0 : boolean;
  signal type_cast_2611_inst_req_1 : boolean;
  signal ptr_deref_2403_load_0_req_0 : boolean;
  signal ptr_deref_2403_load_0_ack_0 : boolean;
  signal type_cast_2611_inst_req_0 : boolean;
  signal ptr_deref_2403_load_0_req_1 : boolean;
  signal ptr_deref_2421_load_0_req_1 : boolean;
  signal ptr_deref_2403_load_0_ack_1 : boolean;
  signal ptr_deref_2421_load_0_ack_1 : boolean;
  signal ptr_deref_2421_load_0_req_0 : boolean;
  signal ptr_deref_2421_load_0_ack_0 : boolean;
  signal type_cast_2611_inst_ack_1 : boolean;
  signal phi_stmt_2605_req_1 : boolean;
  signal RPIPE_Block3_start_2390_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2390_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2390_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2390_inst_ack_1 : boolean;
  signal ptr_deref_2439_load_0_req_0 : boolean;
  signal ptr_deref_2439_load_0_ack_0 : boolean;
  signal ptr_deref_2439_load_0_req_1 : boolean;
  signal ptr_deref_2439_load_0_ack_1 : boolean;
  signal ptr_deref_2449_load_0_req_0 : boolean;
  signal ptr_deref_2449_load_0_ack_0 : boolean;
  signal ptr_deref_2449_load_0_req_1 : boolean;
  signal ptr_deref_2449_load_0_ack_1 : boolean;
  signal ptr_deref_2461_load_0_req_0 : boolean;
  signal ptr_deref_2461_load_0_ack_0 : boolean;
  signal ptr_deref_2461_load_0_req_1 : boolean;
  signal ptr_deref_2461_load_0_ack_1 : boolean;
  signal LOAD_padding_2464_load_0_req_0 : boolean;
  signal LOAD_padding_2464_load_0_ack_0 : boolean;
  signal LOAD_padding_2464_load_0_req_1 : boolean;
  signal LOAD_padding_2464_load_0_ack_1 : boolean;
  signal ptr_deref_2474_load_0_req_0 : boolean;
  signal ptr_deref_2474_load_0_ack_0 : boolean;
  signal ptr_deref_2474_load_0_req_1 : boolean;
  signal ptr_deref_2474_load_0_ack_1 : boolean;
  signal ptr_deref_2486_load_0_req_0 : boolean;
  signal ptr_deref_2486_load_0_ack_0 : boolean;
  signal ptr_deref_2486_load_0_req_1 : boolean;
  signal ptr_deref_2486_load_0_ack_1 : boolean;
  signal ptr_deref_2498_load_0_req_0 : boolean;
  signal ptr_deref_2498_load_0_ack_0 : boolean;
  signal ptr_deref_2498_load_0_req_1 : boolean;
  signal ptr_deref_2498_load_0_ack_1 : boolean;
  signal ptr_deref_2510_load_0_req_0 : boolean;
  signal ptr_deref_2510_load_0_ack_0 : boolean;
  signal ptr_deref_2510_load_0_req_1 : boolean;
  signal ptr_deref_2510_load_0_ack_1 : boolean;
  signal phi_stmt_2605_req_0 : boolean;
  signal type_cast_2514_inst_req_0 : boolean;
  signal type_cast_2514_inst_ack_0 : boolean;
  signal type_cast_2514_inst_req_1 : boolean;
  signal type_cast_2514_inst_ack_1 : boolean;
  signal type_cast_2631_inst_req_0 : boolean;
  signal type_cast_2631_inst_ack_0 : boolean;
  signal type_cast_2631_inst_req_1 : boolean;
  signal type_cast_2631_inst_ack_1 : boolean;
  signal array_obj_ref_2643_index_offset_req_0 : boolean;
  signal array_obj_ref_2643_index_offset_ack_0 : boolean;
  signal array_obj_ref_2643_index_offset_req_1 : boolean;
  signal array_obj_ref_2643_index_offset_ack_1 : boolean;
  signal addr_of_2644_final_reg_req_0 : boolean;
  signal addr_of_2644_final_reg_ack_0 : boolean;
  signal addr_of_2644_final_reg_req_1 : boolean;
  signal addr_of_2644_final_reg_ack_1 : boolean;
  signal ptr_deref_2648_load_0_req_0 : boolean;
  signal ptr_deref_2648_load_0_ack_0 : boolean;
  signal ptr_deref_2648_load_0_req_1 : boolean;
  signal ptr_deref_2648_load_0_ack_1 : boolean;
  signal type_cast_2652_inst_req_0 : boolean;
  signal type_cast_2652_inst_ack_0 : boolean;
  signal type_cast_2652_inst_req_1 : boolean;
  signal type_cast_2652_inst_ack_1 : boolean;
  signal array_obj_ref_2664_index_offset_req_0 : boolean;
  signal array_obj_ref_2664_index_offset_ack_0 : boolean;
  signal array_obj_ref_2664_index_offset_req_1 : boolean;
  signal array_obj_ref_2664_index_offset_ack_1 : boolean;
  signal addr_of_2665_final_reg_req_0 : boolean;
  signal addr_of_2665_final_reg_ack_0 : boolean;
  signal addr_of_2665_final_reg_req_1 : boolean;
  signal addr_of_2665_final_reg_ack_1 : boolean;
  signal ptr_deref_2668_store_0_req_0 : boolean;
  signal ptr_deref_2668_store_0_ack_0 : boolean;
  signal ptr_deref_2668_store_0_req_1 : boolean;
  signal ptr_deref_2668_store_0_ack_1 : boolean;
  signal type_cast_2673_inst_req_0 : boolean;
  signal type_cast_2673_inst_ack_0 : boolean;
  signal type_cast_2673_inst_req_1 : boolean;
  signal type_cast_2673_inst_ack_1 : boolean;
  signal if_stmt_2686_branch_req_0 : boolean;
  signal if_stmt_2686_branch_ack_1 : boolean;
  signal if_stmt_2686_branch_ack_0 : boolean;
  signal if_stmt_2741_branch_req_0 : boolean;
  signal if_stmt_2741_branch_ack_1 : boolean;
  signal if_stmt_2741_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2749_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2749_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2749_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2749_inst_ack_1 : boolean;
  signal type_cast_2545_inst_req_0 : boolean;
  signal type_cast_2545_inst_ack_0 : boolean;
  signal type_cast_2545_inst_req_1 : boolean;
  signal type_cast_2545_inst_ack_1 : boolean;
  signal phi_stmt_2540_req_1 : boolean;
  signal type_cast_2551_inst_req_0 : boolean;
  signal type_cast_2551_inst_ack_0 : boolean;
  signal type_cast_2551_inst_req_1 : boolean;
  signal type_cast_2551_inst_ack_1 : boolean;
  signal phi_stmt_2546_req_1 : boolean;
  signal type_cast_2543_inst_req_0 : boolean;
  signal type_cast_2543_inst_ack_0 : boolean;
  signal type_cast_2543_inst_req_1 : boolean;
  signal type_cast_2543_inst_ack_1 : boolean;
  signal phi_stmt_2540_req_0 : boolean;
  signal type_cast_2549_inst_req_0 : boolean;
  signal type_cast_2549_inst_ack_0 : boolean;
  signal type_cast_2549_inst_req_1 : boolean;
  signal type_cast_2549_inst_ack_1 : boolean;
  signal phi_stmt_2546_req_0 : boolean;
  signal phi_stmt_2540_ack_0 : boolean;
  signal phi_stmt_2546_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7032_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7032_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7032_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7032_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7032: Block -- control-path 
    signal convTransposeD_CP_7032_elements: BooleanArray(75 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7032_elements(0) <= convTransposeD_CP_7032_start;
    convTransposeD_CP_7032_symbol <= convTransposeD_CP_7032_elements(51);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2388/$entry
      -- CP-element group 0: 	 branch_block_stmt_2388/branch_block_stmt_2388__entry__
      -- CP-element group 0: 	 branch_block_stmt_2388/assign_stmt_2391__entry__
      -- CP-element group 0: 	 branch_block_stmt_2388/assign_stmt_2391/$entry
      -- CP-element group 0: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Sample/rr
      -- 
    rr_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(0), ack => RPIPE_Block3_start_2390_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Update/cr
      -- 
    ra_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2390_inst_ack_0, ack => convTransposeD_CP_7032_elements(1)); -- 
    cr_7085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(1), ack => RPIPE_Block3_start_2390_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2:  members (256) 
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2391__exit__
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537__entry__
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2391/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2391/RPIPE_Block3_start_2390_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Update/cr
      -- 
    ca_7086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2390_inst_ack_1, ack => convTransposeD_CP_7032_elements(2)); -- 
    rr_7122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2403_load_0_req_0); -- 
    cr_7133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2403_load_0_req_1); -- 
    cr_7183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2421_load_0_req_1); -- 
    rr_7172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2421_load_0_req_0); -- 
    rr_7222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2439_load_0_req_0); -- 
    cr_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2439_load_0_req_1); -- 
    rr_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2449_load_0_req_0); -- 
    cr_7283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2449_load_0_req_1); -- 
    rr_7322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2461_load_0_req_0); -- 
    cr_7333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2461_load_0_req_1); -- 
    rr_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => LOAD_padding_2464_load_0_req_0); -- 
    cr_7366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => LOAD_padding_2464_load_0_req_1); -- 
    rr_7405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2474_load_0_req_0); -- 
    cr_7416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2474_load_0_req_1); -- 
    rr_7455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2486_load_0_req_0); -- 
    cr_7466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2486_load_0_req_1); -- 
    rr_7505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2498_load_0_req_0); -- 
    cr_7516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2498_load_0_req_1); -- 
    rr_7555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2510_load_0_req_0); -- 
    cr_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => ptr_deref_2510_load_0_req_1); -- 
    cr_7585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(2), ack => type_cast_2514_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_sample_completed_
      -- 
    ra_7123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2403_load_0_ack_0, ack => convTransposeD_CP_7032_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	25 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/ptr_deref_2403_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/ptr_deref_2403_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/ptr_deref_2403_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/ptr_deref_2403_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2403_update_completed_
      -- 
    ca_7134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2403_load_0_ack_1, ack => convTransposeD_CP_7032_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Sample/word_access_start/word_0/ra
      -- 
    ra_7173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2421_load_0_ack_0, ack => convTransposeD_CP_7032_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	25 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/ptr_deref_2421_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/ptr_deref_2421_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/ptr_deref_2421_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/ptr_deref_2421_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2421_Update/word_access_complete/word_0/ca
      -- 
    ca_7184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2421_load_0_ack_1, ack => convTransposeD_CP_7032_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Sample/word_access_start/word_0/ra
      -- 
    ra_7223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2439_load_0_ack_0, ack => convTransposeD_CP_7032_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/ptr_deref_2439_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/ptr_deref_2439_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/ptr_deref_2439_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2439_Update/ptr_deref_2439_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Sample/rr
      -- 
    ca_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2439_load_0_ack_1, ack => convTransposeD_CP_7032_elements(8)); -- 
    rr_7580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(8), ack => type_cast_2514_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Sample/word_access_start/word_0/ra
      -- 
    ra_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2449_load_0_ack_0, ack => convTransposeD_CP_7032_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/ptr_deref_2449_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/ptr_deref_2449_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/ptr_deref_2449_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2449_Update/ptr_deref_2449_Merge/merge_ack
      -- 
    ca_7284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2449_load_0_ack_1, ack => convTransposeD_CP_7032_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Sample/word_access_start/word_0/ra
      -- 
    ra_7323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2461_load_0_ack_0, ack => convTransposeD_CP_7032_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	25 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/ptr_deref_2461_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/ptr_deref_2461_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/ptr_deref_2461_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2461_Update/ptr_deref_2461_Merge/merge_ack
      -- 
    ca_7334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2461_load_0_ack_1, ack => convTransposeD_CP_7032_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Sample/word_access_start/word_0/ra
      -- 
    ra_7356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2464_load_0_ack_0, ack => convTransposeD_CP_7032_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	25 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/LOAD_padding_2464_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/LOAD_padding_2464_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/LOAD_padding_2464_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/LOAD_padding_2464_Update/LOAD_padding_2464_Merge/merge_ack
      -- 
    ca_7367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2464_load_0_ack_1, ack => convTransposeD_CP_7032_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Sample/word_access_start/word_0/ra
      -- 
    ra_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2474_load_0_ack_0, ack => convTransposeD_CP_7032_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	25 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/ptr_deref_2474_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/ptr_deref_2474_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/ptr_deref_2474_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2474_Update/ptr_deref_2474_Merge/merge_ack
      -- 
    ca_7417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2474_load_0_ack_1, ack => convTransposeD_CP_7032_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Sample/word_access_start/word_0/ra
      -- 
    ra_7456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2486_load_0_ack_0, ack => convTransposeD_CP_7032_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/ptr_deref_2486_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/ptr_deref_2486_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/ptr_deref_2486_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2486_Update/ptr_deref_2486_Merge/merge_ack
      -- 
    ca_7467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2486_load_0_ack_1, ack => convTransposeD_CP_7032_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Sample/word_access_start/word_0/ra
      -- 
    ra_7506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2498_load_0_ack_0, ack => convTransposeD_CP_7032_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/ptr_deref_2498_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/ptr_deref_2498_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/ptr_deref_2498_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2498_Update/ptr_deref_2498_Merge/merge_ack
      -- 
    ca_7517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2498_load_0_ack_1, ack => convTransposeD_CP_7032_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Sample/word_access_start/word_0/ra
      -- 
    ra_7556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2510_load_0_ack_0, ack => convTransposeD_CP_7032_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/ptr_deref_2510_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/ptr_deref_2510_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/ptr_deref_2510_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/ptr_deref_2510_Update/ptr_deref_2510_Merge/merge_ack
      -- 
    ca_7567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2510_load_0_ack_1, ack => convTransposeD_CP_7032_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Sample/ra
      -- 
    ra_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2514_inst_ack_0, ack => convTransposeD_CP_7032_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/type_cast_2514_Update/ca
      -- 
    ca_7586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2514_inst_ack_1, ack => convTransposeD_CP_7032_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  place  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: 	18 
    -- CP-element group 25: 	22 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	12 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	14 
    -- CP-element group 25: 	4 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	55 
    -- CP-element group 25: 	56 
    -- CP-element group 25: 	52 
    -- CP-element group 25: 	53 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537__exit__
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter
      -- CP-element group 25: 	 branch_block_stmt_2388/assign_stmt_2400_to_assign_stmt_2537/$exit
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Update/cr
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Update/cr
      -- 
    rr_7906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(25), ack => type_cast_2545_inst_req_0); -- 
    cr_7911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(25), ack => type_cast_2545_inst_req_1); -- 
    rr_7929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(25), ack => type_cast_2551_inst_req_0); -- 
    cr_7934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(25), ack => type_cast_2551_inst_req_1); -- 
    convTransposeD_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(24) & convTransposeD_CP_7032_elements(18) & convTransposeD_CP_7032_elements(22) & convTransposeD_CP_7032_elements(20) & convTransposeD_CP_7032_elements(12) & convTransposeD_CP_7032_elements(16) & convTransposeD_CP_7032_elements(14) & convTransposeD_CP_7032_elements(4) & convTransposeD_CP_7032_elements(6) & convTransposeD_CP_7032_elements(10);
      gj_convTransposeD_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	75 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Sample/ra
      -- 
    ra_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_0, ack => convTransposeD_CP_7032_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	75 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (16) 
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Sample/req
      -- 
    ca_7606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_1, ack => convTransposeD_CP_7032_elements(27)); -- 
    req_7631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(27), ack => array_obj_ref_2643_index_offset_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	45 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_sample_complete
      -- CP-element group 28: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Sample/ack
      -- 
    ack_7632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2643_index_offset_ack_0, ack => convTransposeD_CP_7032_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	75 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (11) 
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_root_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_offset_calculated
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_base_plus_offset/$entry
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_base_plus_offset/$exit
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_base_plus_offset/sum_rename_req
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_base_plus_offset/sum_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_request/$entry
      -- CP-element group 29: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_request/req
      -- 
    ack_7637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2643_index_offset_ack_1, ack => convTransposeD_CP_7032_elements(29)); -- 
    req_7646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(29), ack => addr_of_2644_final_reg_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_request/$exit
      -- CP-element group 30: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_request/ack
      -- 
    ack_7647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2644_final_reg_ack_0, ack => convTransposeD_CP_7032_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	75 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (24) 
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_complete/ack
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_address_resized
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_addr_resize/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_addr_resize/$exit
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_addr_resize/base_resize_req
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_addr_resize/base_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_word_addrgen/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_word_addrgen/$exit
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_word_addrgen/root_register_req
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_word_addrgen/root_register_ack
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/word_0/rr
      -- 
    ack_7652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2644_final_reg_ack_1, ack => convTransposeD_CP_7032_elements(31)); -- 
    rr_7685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(31), ack => ptr_deref_2648_load_0_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Sample/word_access_start/word_0/ra
      -- 
    ra_7686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_load_0_ack_0, ack => convTransposeD_CP_7032_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	40 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/word_0/ca
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/ptr_deref_2648_Merge/$entry
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/ptr_deref_2648_Merge/$exit
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/ptr_deref_2648_Merge/merge_req
      -- CP-element group 33: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/ptr_deref_2648_Merge/merge_ack
      -- 
    ca_7697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2648_load_0_ack_1, ack => convTransposeD_CP_7032_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	75 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Sample/ra
      -- 
    ra_7711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2652_inst_ack_0, ack => convTransposeD_CP_7032_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	75 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Sample/req
      -- 
    ca_7716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2652_inst_ack_1, ack => convTransposeD_CP_7032_elements(35)); -- 
    req_7741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(35), ack => array_obj_ref_2664_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Sample/ack
      -- 
    ack_7742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2664_index_offset_ack_0, ack => convTransposeD_CP_7032_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	75 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_request/req
      -- 
    ack_7747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2664_index_offset_ack_1, ack => convTransposeD_CP_7032_elements(37)); -- 
    req_7756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(37), ack => addr_of_2665_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_request/ack
      -- 
    ack_7757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2665_final_reg_ack_0, ack => convTransposeD_CP_7032_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	75 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (19) 
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_word_addrgen/root_register_ack
      -- 
    ack_7762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2665_final_reg_ack_1, ack => convTransposeD_CP_7032_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: 	33 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/ptr_deref_2668_Split/$entry
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/ptr_deref_2668_Split/$exit
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/ptr_deref_2668_Split/split_req
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/ptr_deref_2668_Split/split_ack
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/$entry
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/word_0/rr
      -- 
    rr_7800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(40), ack => ptr_deref_2668_store_0_req_0); -- 
    convTransposeD_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(39) & convTransposeD_CP_7032_elements(33);
      gj_convTransposeD_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/$exit
      -- CP-element group 41: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Sample/word_access_start/word_0/ra
      -- 
    ra_7801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2668_store_0_ack_0, ack => convTransposeD_CP_7032_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	75 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/word_0/ca
      -- 
    ca_7812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2668_store_0_ack_1, ack => convTransposeD_CP_7032_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	75 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Sample/ra
      -- 
    ra_7821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2673_inst_ack_0, ack => convTransposeD_CP_7032_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	75 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Update/ca
      -- 
    ca_7826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2673_inst_ack_1, ack => convTransposeD_CP_7032_elements(44)); -- 
    -- CP-element group 45:  branch  join  transition  place  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	28 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (10) 
      -- CP-element group 45: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685__exit__
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686__entry__
      -- CP-element group 45: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/$exit
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_dead_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_eval_test/$entry
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_eval_test/$exit
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_eval_test/branch_req
      -- CP-element group 45: 	 branch_block_stmt_2388/R_cmp_2687_place
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_if_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_2388/if_stmt_2686_else_link/$entry
      -- 
    branch_req_7834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(45), ack => if_stmt_2686_branch_req_0); -- 
    convTransposeD_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(36) & convTransposeD_CP_7032_elements(44) & convTransposeD_CP_7032_elements(28) & convTransposeD_CP_7032_elements(42);
      gj_convTransposeD_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	70 
    -- CP-element group 46: 	71 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2388/merge_stmt_2692_PhiAck/dummy
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Update/cr
      -- CP-element group 46: 	 branch_block_stmt_2388/merge_stmt_2692_PhiAck/$exit
      -- CP-element group 46: 	 branch_block_stmt_2388/merge_stmt_2692_PhiAck/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_2388/merge_stmt_2692_PhiReqMerge
      -- CP-element group 46: 	 branch_block_stmt_2388/merge_stmt_2692__exit__
      -- CP-element group 46: 	 branch_block_stmt_2388/assign_stmt_2698__entry__
      -- CP-element group 46: 	 branch_block_stmt_2388/assign_stmt_2698__exit__
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 46: 	 branch_block_stmt_2388/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/if_stmt_2686_if_link/$exit
      -- CP-element group 46: 	 branch_block_stmt_2388/if_stmt_2686_if_link/if_choice_transition
      -- CP-element group 46: 	 branch_block_stmt_2388/whilex_xbody_ifx_xthen
      -- CP-element group 46: 	 branch_block_stmt_2388/assign_stmt_2698/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/assign_stmt_2698/$exit
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/$entry
      -- CP-element group 46: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/$entry
      -- 
    if_choice_transition_7839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2686_branch_ack_1, ack => convTransposeD_CP_7032_elements(46)); -- 
    cr_8015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(46), ack => type_cast_2611_inst_req_1); -- 
    rr_8010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(46), ack => type_cast_2611_inst_req_0); -- 
    -- CP-element group 47:  branch  transition  place  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (22) 
      -- CP-element group 47: 	 branch_block_stmt_2388/merge_stmt_2700_PhiAck/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/merge_stmt_2700_PhiReqMerge
      -- CP-element group 47: 	 branch_block_stmt_2388/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 47: 	 branch_block_stmt_2388/merge_stmt_2700_PhiAck/$exit
      -- CP-element group 47: 	 branch_block_stmt_2388/merge_stmt_2700_PhiAck/dummy
      -- CP-element group 47: 	 branch_block_stmt_2388/merge_stmt_2700__exit__
      -- CP-element group 47: 	 branch_block_stmt_2388/assign_stmt_2706_to_assign_stmt_2740__entry__
      -- CP-element group 47: 	 branch_block_stmt_2388/assign_stmt_2706_to_assign_stmt_2740__exit__
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741__entry__
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2686_else_link/$exit
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2686_else_link/else_choice_transition
      -- CP-element group 47: 	 branch_block_stmt_2388/whilex_xbody_ifx_xelse
      -- CP-element group 47: 	 branch_block_stmt_2388/assign_stmt_2706_to_assign_stmt_2740/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/assign_stmt_2706_to_assign_stmt_2740/$exit
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_2388/R_cmp104_2742_place
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2388/if_stmt_2741_else_link/$entry
      -- 
    else_choice_transition_7843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2686_branch_ack_0, ack => convTransposeD_CP_7032_elements(47)); -- 
    branch_req_7859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(47), ack => if_stmt_2741_branch_req_0); -- 
    -- CP-element group 48:  merge  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (15) 
      -- CP-element group 48: 	 branch_block_stmt_2388/merge_stmt_2747_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_2388/merge_stmt_2747_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_2388/merge_stmt_2747_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_2388/merge_stmt_2747_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_2388/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2388/merge_stmt_2747__exit__
      -- CP-element group 48: 	 branch_block_stmt_2388/assign_stmt_2751__entry__
      -- CP-element group 48: 	 branch_block_stmt_2388/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_2388/if_stmt_2741_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_2388/if_stmt_2741_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_2388/ifx_xelse_whilex_xend
      -- CP-element group 48: 	 branch_block_stmt_2388/assign_stmt_2751/$entry
      -- CP-element group 48: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Sample/req
      -- 
    if_choice_transition_7864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2741_branch_ack_1, ack => convTransposeD_CP_7032_elements(48)); -- 
    req_7881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(48), ack => WPIPE_Block3_done_2749_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	59 
    -- CP-element group 49: 	60 
    -- CP-element group 49: 	62 
    -- CP-element group 49: 	63 
    -- CP-element group 49:  members (20) 
      -- CP-element group 49: 	 branch_block_stmt_2388/if_stmt_2741_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_2388/if_stmt_2741_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Update/cr
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2741_branch_ack_0, ack => convTransposeD_CP_7032_elements(49)); -- 
    rr_7955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(49), ack => type_cast_2543_inst_req_0); -- 
    cr_7960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(49), ack => type_cast_2543_inst_req_1); -- 
    rr_7978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(49), ack => type_cast_2549_inst_req_0); -- 
    cr_7983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(49), ack => type_cast_2549_inst_req_1); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Update/req
      -- 
    ack_7882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2749_inst_ack_0, ack => convTransposeD_CP_7032_elements(50)); -- 
    req_7886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(50), ack => WPIPE_Block3_done_2749_inst_req_1); -- 
    -- CP-element group 51:  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2388/merge_stmt_2753_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_2388/return___PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_2388/return___PhiReq/$exit
      -- CP-element group 51: 	 $exit
      -- CP-element group 51: 	 branch_block_stmt_2388/$exit
      -- CP-element group 51: 	 branch_block_stmt_2388/branch_block_stmt_2388__exit__
      -- CP-element group 51: 	 branch_block_stmt_2388/assign_stmt_2751__exit__
      -- CP-element group 51: 	 branch_block_stmt_2388/return__
      -- CP-element group 51: 	 branch_block_stmt_2388/merge_stmt_2753__exit__
      -- CP-element group 51: 	 branch_block_stmt_2388/merge_stmt_2753_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_2388/merge_stmt_2753_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_2388/merge_stmt_2753_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_2388/assign_stmt_2751/$exit
      -- CP-element group 51: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2388/assign_stmt_2751/WPIPE_Block3_done_2749_Update/ack
      -- 
    ack_7887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2749_inst_ack_1, ack => convTransposeD_CP_7032_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	25 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Sample/ra
      -- 
    ra_7907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_0, ack => convTransposeD_CP_7032_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	25 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/Update/ca
      -- 
    ca_7912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2545_inst_ack_1, ack => convTransposeD_CP_7032_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	58 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/$exit
      -- CP-element group 54: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/$exit
      -- CP-element group 54: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/$exit
      -- CP-element group 54: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2545/SplitProtocol/$exit
      -- CP-element group 54: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_req
      -- 
    phi_stmt_2540_req_7913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2540_req_7913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(54), ack => phi_stmt_2540_req_1); -- 
    convTransposeD_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(52) & convTransposeD_CP_7032_elements(53);
      gj_convTransposeD_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	25 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Sample/ra
      -- 
    ra_7930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2551_inst_ack_0, ack => convTransposeD_CP_7032_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	25 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/Update/ca
      -- 
    ca_7935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2551_inst_ack_1, ack => convTransposeD_CP_7032_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/$exit
      -- CP-element group 57: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/$exit
      -- CP-element group 57: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/$exit
      -- CP-element group 57: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2551/SplitProtocol/$exit
      -- CP-element group 57: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_req
      -- 
    phi_stmt_2546_req_7936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2546_req_7936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(57), ack => phi_stmt_2546_req_1); -- 
    convTransposeD_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(55) & convTransposeD_CP_7032_elements(56);
      gj_convTransposeD_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	54 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2388/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(57) & convTransposeD_CP_7032_elements(54);
      gj_convTransposeD_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	49 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Sample/ra
      -- 
    ra_7956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_0, ack => convTransposeD_CP_7032_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	49 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/Update/ca
      -- 
    ca_7961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_1, ack => convTransposeD_CP_7032_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	65 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/$exit
      -- CP-element group 61: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/$exit
      -- CP-element group 61: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/$exit
      -- CP-element group 61: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_sources/type_cast_2543/SplitProtocol/$exit
      -- CP-element group 61: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2540/phi_stmt_2540_req
      -- 
    phi_stmt_2540_req_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2540_req_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(61), ack => phi_stmt_2540_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(59) & convTransposeD_CP_7032_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	49 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Sample/ra
      -- 
    ra_7979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_0, ack => convTransposeD_CP_7032_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	49 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/Update/ca
      -- 
    ca_7984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_1, ack => convTransposeD_CP_7032_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/$exit
      -- CP-element group 64: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/$exit
      -- CP-element group 64: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/$exit
      -- CP-element group 64: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_sources/type_cast_2549/SplitProtocol/$exit
      -- CP-element group 64: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2546/phi_stmt_2546_req
      -- 
    phi_stmt_2546_req_7985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2546_req_7985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(64), ack => phi_stmt_2546_req_0); -- 
    convTransposeD_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(62) & convTransposeD_CP_7032_elements(63);
      gj_convTransposeD_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	61 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2388/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(61) & convTransposeD_CP_7032_elements(64);
      gj_convTransposeD_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  fork  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	58 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_2388/merge_stmt_2539_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_2388/merge_stmt_2539_PhiAck/$entry
      -- 
    convTransposeD_CP_7032_elements(66) <= OrReduce(convTransposeD_CP_7032_elements(58) & convTransposeD_CP_7032_elements(65));
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2388/merge_stmt_2539_PhiAck/phi_stmt_2540_ack
      -- 
    phi_stmt_2540_ack_7990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2540_ack_0, ack => convTransposeD_CP_7032_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2388/merge_stmt_2539_PhiAck/phi_stmt_2546_ack
      -- 
    phi_stmt_2546_ack_7991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2546_ack_0, ack => convTransposeD_CP_7032_elements(68)); -- 
    -- CP-element group 69:  join  transition  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2388/merge_stmt_2539__exit__
      -- CP-element group 69: 	 branch_block_stmt_2388/assign_stmt_2557_to_assign_stmt_2602__entry__
      -- CP-element group 69: 	 branch_block_stmt_2388/assign_stmt_2557_to_assign_stmt_2602__exit__
      -- CP-element group 69: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 69: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/$entry
      -- CP-element group 69: 	 branch_block_stmt_2388/assign_stmt_2557_to_assign_stmt_2602/$entry
      -- CP-element group 69: 	 branch_block_stmt_2388/assign_stmt_2557_to_assign_stmt_2602/$exit
      -- CP-element group 69: 	 branch_block_stmt_2388/merge_stmt_2539_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(67) & convTransposeD_CP_7032_elements(68);
      gj_convTransposeD_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	46 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Sample/ra
      -- 
    ra_8011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2611_inst_ack_0, ack => convTransposeD_CP_7032_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	46 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/Update/ca
      -- 
    ca_8016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2611_inst_ack_1, ack => convTransposeD_CP_7032_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_req
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/SplitProtocol/$exit
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/$exit
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_2388/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2611/$exit
      -- 
    phi_stmt_2605_req_8017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2605_req_8017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(72), ack => phi_stmt_2605_req_1); -- 
    convTransposeD_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7032_elements(70) & convTransposeD_CP_7032_elements(71);
      gj_convTransposeD_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7032_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 73: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_req
      -- CP-element group 73: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/type_cast_2609_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/phi_stmt_2605_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2388/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2605/$exit
      -- 
    phi_stmt_2605_req_8028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2605_req_8028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(73), ack => phi_stmt_2605_req_0); -- 
    -- Element group convTransposeD_CP_7032_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeD_CP_7032_elements(69), ack => convTransposeD_CP_7032_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  merge  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2388/merge_stmt_2604_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2388/merge_stmt_2604_PhiReqMerge
      -- 
    convTransposeD_CP_7032_elements(74) <= OrReduce(convTransposeD_CP_7032_elements(72) & convTransposeD_CP_7032_elements(73));
    -- CP-element group 75:  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	29 
    -- CP-element group 75: 	39 
    -- CP-element group 75: 	44 
    -- CP-element group 75: 	31 
    -- CP-element group 75: 	26 
    -- CP-element group 75: 	33 
    -- CP-element group 75: 	37 
    -- CP-element group 75: 	34 
    -- CP-element group 75: 	35 
    -- CP-element group 75: 	27 
    -- CP-element group 75: 	42 
    -- CP-element group 75: 	43 
    -- CP-element group 75:  members (45) 
      -- CP-element group 75: 	 branch_block_stmt_2388/merge_stmt_2604_PhiAck/phi_stmt_2605_ack
      -- CP-element group 75: 	 branch_block_stmt_2388/merge_stmt_2604_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2388/merge_stmt_2604__exit__
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685__entry__
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2631_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_update_start
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2643_final_index_sum_regn_Update/req
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2644_complete/req
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2648_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2652_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_update_start
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/array_obj_ref_2664_final_index_sum_regn_Update/req
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/addr_of_2665_complete/req
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/ptr_deref_2668_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2388/assign_stmt_2618_to_assign_stmt_2685/type_cast_2673_Update/cr
      -- 
    phi_stmt_2605_ack_8033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2605_ack_0, ack => convTransposeD_CP_7032_elements(75)); -- 
    rr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2631_inst_req_0); -- 
    cr_7605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2631_inst_req_1); -- 
    req_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => array_obj_ref_2643_index_offset_req_1); -- 
    req_7651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => addr_of_2644_final_reg_req_1); -- 
    cr_7696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => ptr_deref_2648_load_0_req_1); -- 
    rr_7710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2652_inst_req_0); -- 
    cr_7715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2652_inst_req_1); -- 
    req_7746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => array_obj_ref_2664_index_offset_req_1); -- 
    req_7761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => addr_of_2665_final_reg_req_1); -- 
    cr_7811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => ptr_deref_2668_store_0_req_1); -- 
    rr_7820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2673_inst_req_0); -- 
    cr_7825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7032_elements(75), ack => type_cast_2673_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_2464_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2464_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr118_2642_resized : std_logic_vector(13 downto 0);
    signal R_shr118_2642_scaled : std_logic_vector(13 downto 0);
    signal R_shr72120_2663_resized : std_logic_vector(13 downto 0);
    signal R_shr72120_2663_scaled : std_logic_vector(13 downto 0);
    signal add25_2623 : std_logic_vector(15 downto 0);
    signal add65_2628 : std_logic_vector(15 downto 0);
    signal add78_2680 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2643_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2643_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2643_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2643_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2643_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2643_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2664_root_address : std_logic_vector(13 downto 0);
    signal arrayidx74_2666 : std_logic_vector(31 downto 0);
    signal arrayidx_2645 : std_logic_vector(31 downto 0);
    signal call_2391 : std_logic_vector(15 downto 0);
    signal cmp104_2740 : std_logic_vector(0 downto 0);
    signal cmp91_2711 : std_logic_vector(0 downto 0);
    signal cmp_2685 : std_logic_vector(0 downto 0);
    signal conv68_2632 : std_logic_vector(63 downto 0);
    signal conv71_2653 : std_logic_vector(63 downto 0);
    signal conv77_2674 : std_logic_vector(31 downto 0);
    signal conv80_2515 : std_logic_vector(31 downto 0);
    signal div5_2428 : std_logic_vector(15 downto 0);
    signal div98_2723 : std_logic_vector(15 downto 0);
    signal div_2410 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2507 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2400 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2418 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2436 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2446 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2458 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2471 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2483 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2495 : std_logic_vector(31 downto 0);
    signal inc95_2717 : std_logic_vector(15 downto 0);
    signal inc_2706 : std_logic_vector(15 downto 0);
    signal indvar_2605 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2698 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2735 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2546 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2540 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2729 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2618 : std_logic_vector(15 downto 0);
    signal ptr_deref_2403_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2403_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2421_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2421_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2439_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2439_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2439_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2439_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2439_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2449_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2449_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2449_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2449_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2449_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2461_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2461_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2461_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2461_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2461_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2474_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2474_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2474_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2474_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2474_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2486_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2486_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2486_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2498_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2498_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2510_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2510_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2510_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2510_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2510_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2648_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2648_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2648_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2648_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2648_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2668_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2668_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2668_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2668_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2668_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2668_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr118_2638 : std_logic_vector(63 downto 0);
    signal shr72120_2659 : std_logic_vector(63 downto 0);
    signal tmp10_2582 : std_logic_vector(15 downto 0);
    signal tmp11_2587 : std_logic_vector(15 downto 0);
    signal tmp12_2592 : std_logic_vector(15 downto 0);
    signal tmp134_2557 : std_logic_vector(15 downto 0);
    signal tmp135_2562 : std_logic_vector(15 downto 0);
    signal tmp136_2567 : std_logic_vector(15 downto 0);
    signal tmp13_2597 : std_logic_vector(15 downto 0);
    signal tmp14_2602 : std_logic_vector(15 downto 0);
    signal tmp16_2440 : std_logic_vector(15 downto 0);
    signal tmp29_2450 : std_logic_vector(15 downto 0);
    signal tmp32_2462 : std_logic_vector(15 downto 0);
    signal tmp35_2465 : std_logic_vector(15 downto 0);
    signal tmp3_2422 : std_logic_vector(15 downto 0);
    signal tmp41_2475 : std_logic_vector(15 downto 0);
    signal tmp44_2487 : std_logic_vector(15 downto 0);
    signal tmp4_2521 : std_logic_vector(15 downto 0);
    signal tmp54_2499 : std_logic_vector(15 downto 0);
    signal tmp58_2511 : std_logic_vector(15 downto 0);
    signal tmp5_2526 : std_logic_vector(15 downto 0);
    signal tmp69_2649 : std_logic_vector(63 downto 0);
    signal tmp6_2572 : std_logic_vector(15 downto 0);
    signal tmp7_2577 : std_logic_vector(15 downto 0);
    signal tmp8_2532 : std_logic_vector(15 downto 0);
    signal tmp9_2537 : std_logic_vector(15 downto 0);
    signal tmp_2404 : std_logic_vector(15 downto 0);
    signal type_cast_2408_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2426_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2519_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2530_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2543_wire : std_logic_vector(15 downto 0);
    signal type_cast_2545_wire : std_logic_vector(15 downto 0);
    signal type_cast_2549_wire : std_logic_vector(15 downto 0);
    signal type_cast_2551_wire : std_logic_vector(15 downto 0);
    signal type_cast_2609_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2611_wire : std_logic_vector(15 downto 0);
    signal type_cast_2616_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2636_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2657_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2678_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2696_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2704_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2715_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_2464_word_address_0 <= "0";
    array_obj_ref_2643_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2643_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2643_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2643_resized_base_address <= "00000000000000";
    array_obj_ref_2664_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2664_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2664_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2664_resized_base_address <= "00000000000000";
    iNsTr_10_2507 <= "00000000000000000000000000000100";
    iNsTr_2_2400 <= "00000000000000000000000000000011";
    iNsTr_3_2418 <= "00000000000000000000000000000100";
    iNsTr_4_2436 <= "00000000000000000000000000000101";
    iNsTr_5_2446 <= "00000000000000000000000000000000";
    iNsTr_6_2458 <= "00000000000000000000000000000100";
    iNsTr_7_2471 <= "00000000000000000000000000000001";
    iNsTr_8_2483 <= "00000000000000000000000000000101";
    iNsTr_9_2495 <= "00000000000000000000000000000101";
    ptr_deref_2403_word_offset_0 <= "0000000";
    ptr_deref_2421_word_offset_0 <= "0000000";
    ptr_deref_2439_word_offset_0 <= "0000000";
    ptr_deref_2449_word_offset_0 <= "0";
    ptr_deref_2461_word_offset_0 <= "0000000";
    ptr_deref_2474_word_offset_0 <= "0";
    ptr_deref_2486_word_offset_0 <= "0000000";
    ptr_deref_2498_word_offset_0 <= "0000000";
    ptr_deref_2510_word_offset_0 <= "0000000";
    ptr_deref_2648_word_offset_0 <= "00000000000000";
    ptr_deref_2668_word_offset_0 <= "00000000000000";
    type_cast_2408_wire_constant <= "0000000000000001";
    type_cast_2426_wire_constant <= "0000000000000001";
    type_cast_2519_wire_constant <= "1111111111111111";
    type_cast_2530_wire_constant <= "1111111111111111";
    type_cast_2609_wire_constant <= "0000000000000000";
    type_cast_2616_wire_constant <= "0000000000000100";
    type_cast_2636_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2657_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2678_wire_constant <= "00000000000000000000000000000100";
    type_cast_2696_wire_constant <= "0000000000000001";
    type_cast_2704_wire_constant <= "0000000000000001";
    type_cast_2715_wire_constant <= "0000000000000001";
    type_cast_2721_wire_constant <= "0000000000000001";
    phi_stmt_2540: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2543_wire & type_cast_2545_wire;
      req <= phi_stmt_2540_req_0 & phi_stmt_2540_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2540",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2540_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2540,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2540
    phi_stmt_2546: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2549_wire & type_cast_2551_wire;
      req <= phi_stmt_2546_req_0 & phi_stmt_2546_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2546",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2546_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2546,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2546
    phi_stmt_2605: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2609_wire_constant & type_cast_2611_wire;
      req <= phi_stmt_2605_req_0 & phi_stmt_2605_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2605",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2605_ack_0,
          idata => idata,
          odata => indvar_2605,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2605
    -- flow-through select operator MUX_2728_inst
    input_dim1x_x2_2729 <= div98_2723 when (cmp91_2711(0) /=  '0') else inc_2706;
    -- flow-through select operator MUX_2734_inst
    input_dim0x_x0_2735 <= inc95_2717 when (cmp91_2711(0) /=  '0') else input_dim0x_x2x_xph_2546;
    addr_of_2644_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2644_final_reg_req_0;
      addr_of_2644_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2644_final_reg_req_1;
      addr_of_2644_final_reg_ack_1<= rack(0);
      addr_of_2644_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2644_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2643_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2665_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2665_final_reg_req_0;
      addr_of_2665_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2665_final_reg_req_1;
      addr_of_2665_final_reg_ack_1<= rack(0);
      addr_of_2665_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2665_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2664_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx74_2666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2514_inst_req_0;
      type_cast_2514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2514_inst_req_1;
      type_cast_2514_inst_ack_1<= rack(0);
      type_cast_2514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2543_inst_req_0;
      type_cast_2543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2543_inst_req_1;
      type_cast_2543_inst_ack_1<= rack(0);
      type_cast_2543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2543_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2545_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2545_inst_req_0;
      type_cast_2545_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2545_inst_req_1;
      type_cast_2545_inst_ack_1<= rack(0);
      type_cast_2545_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2545_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div5_2428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2545_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2549_inst_req_0;
      type_cast_2549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2549_inst_req_1;
      type_cast_2549_inst_ack_1<= rack(0);
      type_cast_2549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2549_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2551_inst_req_0;
      type_cast_2551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2551_inst_req_1;
      type_cast_2551_inst_ack_1<= rack(0);
      type_cast_2551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2551_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2611_inst_req_0;
      type_cast_2611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2611_inst_req_1;
      type_cast_2611_inst_ack_1<= rack(0);
      type_cast_2611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2611_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2631_inst_req_0;
      type_cast_2631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2631_inst_req_1;
      type_cast_2631_inst_ack_1<= rack(0);
      type_cast_2631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add25_2623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2652_inst_req_0;
      type_cast_2652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2652_inst_req_1;
      type_cast_2652_inst_ack_1<= rack(0);
      type_cast_2652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add65_2628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_2653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2673_inst_req_0;
      type_cast_2673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2673_inst_req_1;
      type_cast_2673_inst_ack_1<= rack(0);
      type_cast_2673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_2674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2464_gather_scatter
    process(LOAD_padding_2464_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2464_data_0;
      ov(15 downto 0) := iv;
      tmp35_2465 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2643_index_1_rename
    process(R_shr118_2642_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr118_2642_resized;
      ov(13 downto 0) := iv;
      R_shr118_2642_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2643_index_1_resize
    process(shr118_2638) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr118_2638;
      ov := iv(13 downto 0);
      R_shr118_2642_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2643_root_address_inst
    process(array_obj_ref_2643_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2643_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2643_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2664_index_1_rename
    process(R_shr72120_2663_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr72120_2663_resized;
      ov(13 downto 0) := iv;
      R_shr72120_2663_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2664_index_1_resize
    process(shr72120_2659) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr72120_2659;
      ov := iv(13 downto 0);
      R_shr72120_2663_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2664_root_address_inst
    process(array_obj_ref_2664_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2664_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2664_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_addr_0
    process(ptr_deref_2403_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2403_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_base_resize
    process(iNsTr_2_2400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2400;
      ov := iv(6 downto 0);
      ptr_deref_2403_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_gather_scatter
    process(ptr_deref_2403_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_data_0;
      ov(15 downto 0) := iv;
      tmp_2404 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_root_address_inst
    process(ptr_deref_2403_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2403_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_addr_0
    process(ptr_deref_2421_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2421_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_base_resize
    process(iNsTr_3_2418) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2418;
      ov := iv(6 downto 0);
      ptr_deref_2421_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_gather_scatter
    process(ptr_deref_2421_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_data_0;
      ov(15 downto 0) := iv;
      tmp3_2422 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2421_root_address_inst
    process(ptr_deref_2421_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2421_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2421_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2439_addr_0
    process(ptr_deref_2439_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2439_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2439_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2439_base_resize
    process(iNsTr_4_2436) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2436;
      ov := iv(6 downto 0);
      ptr_deref_2439_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2439_gather_scatter
    process(ptr_deref_2439_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2439_data_0;
      ov(15 downto 0) := iv;
      tmp16_2440 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2439_root_address_inst
    process(ptr_deref_2439_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2439_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2439_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_addr_0
    process(ptr_deref_2449_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2449_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_base_resize
    process(iNsTr_5_2446) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2446;
      ov := iv(0 downto 0);
      ptr_deref_2449_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_gather_scatter
    process(ptr_deref_2449_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_data_0;
      ov(15 downto 0) := iv;
      tmp29_2450 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2449_root_address_inst
    process(ptr_deref_2449_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2449_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2449_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2461_addr_0
    process(ptr_deref_2461_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2461_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2461_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2461_base_resize
    process(iNsTr_6_2458) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2458;
      ov := iv(6 downto 0);
      ptr_deref_2461_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2461_gather_scatter
    process(ptr_deref_2461_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2461_data_0;
      ov(15 downto 0) := iv;
      tmp32_2462 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2461_root_address_inst
    process(ptr_deref_2461_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2461_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2461_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2474_addr_0
    process(ptr_deref_2474_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2474_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2474_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2474_base_resize
    process(iNsTr_7_2471) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2471;
      ov := iv(0 downto 0);
      ptr_deref_2474_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2474_gather_scatter
    process(ptr_deref_2474_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2474_data_0;
      ov(15 downto 0) := iv;
      tmp41_2475 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2474_root_address_inst
    process(ptr_deref_2474_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2474_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2474_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_addr_0
    process(ptr_deref_2486_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2486_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_base_resize
    process(iNsTr_8_2483) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2483;
      ov := iv(6 downto 0);
      ptr_deref_2486_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_gather_scatter
    process(ptr_deref_2486_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_data_0;
      ov(15 downto 0) := iv;
      tmp44_2487 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2486_root_address_inst
    process(ptr_deref_2486_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2486_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2486_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_addr_0
    process(ptr_deref_2498_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2498_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_base_resize
    process(iNsTr_9_2495) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2495;
      ov := iv(6 downto 0);
      ptr_deref_2498_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_gather_scatter
    process(ptr_deref_2498_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_data_0;
      ov(15 downto 0) := iv;
      tmp54_2499 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2498_root_address_inst
    process(ptr_deref_2498_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2498_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2498_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2510_addr_0
    process(ptr_deref_2510_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2510_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2510_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2510_base_resize
    process(iNsTr_10_2507) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2507;
      ov := iv(6 downto 0);
      ptr_deref_2510_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2510_gather_scatter
    process(ptr_deref_2510_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2510_data_0;
      ov(15 downto 0) := iv;
      tmp58_2511 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2510_root_address_inst
    process(ptr_deref_2510_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2510_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2510_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2648_addr_0
    process(ptr_deref_2648_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2648_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2648_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2648_base_resize
    process(arrayidx_2645) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2645;
      ov := iv(13 downto 0);
      ptr_deref_2648_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2648_gather_scatter
    process(ptr_deref_2648_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2648_data_0;
      ov(63 downto 0) := iv;
      tmp69_2649 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2648_root_address_inst
    process(ptr_deref_2648_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2648_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2648_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2668_addr_0
    process(ptr_deref_2668_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2668_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2668_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2668_base_resize
    process(arrayidx74_2666) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx74_2666;
      ov := iv(13 downto 0);
      ptr_deref_2668_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2668_gather_scatter
    process(tmp69_2649) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp69_2649;
      ov(63 downto 0) := iv;
      ptr_deref_2668_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2668_root_address_inst
    process(ptr_deref_2668_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2668_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2668_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2686_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2685;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2686_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2686_branch_req_0,
          ack0 => if_stmt_2686_branch_ack_0,
          ack1 => if_stmt_2686_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2741_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp104_2740;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2741_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2741_branch_req_0,
          ack0 => if_stmt_2741_branch_ack_0,
          ack1 => if_stmt_2741_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2520_inst
    process(tmp44_2487) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp44_2487, type_cast_2519_wire_constant, tmp_var);
      tmp4_2521 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2531_inst
    process(tmp32_2462) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp32_2462, type_cast_2530_wire_constant, tmp_var);
      tmp8_2532 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2561_inst
    process(input_dim1x_x1x_xph_2540, tmp134_2557) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2540, tmp134_2557, tmp_var);
      tmp135_2562 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2576_inst
    process(tmp5_2526, tmp6_2572) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2526, tmp6_2572, tmp_var);
      tmp7_2577 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2586_inst
    process(tmp9_2537, tmp10_2582) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_2537, tmp10_2582, tmp_var);
      tmp11_2587 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2596_inst
    process(tmp7_2577, tmp12_2592) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_2577, tmp12_2592, tmp_var);
      tmp13_2597 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2622_inst
    process(tmp136_2567, input_dim2x_x1_2618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp136_2567, input_dim2x_x1_2618, tmp_var);
      add25_2623 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2627_inst
    process(tmp14_2602, input_dim2x_x1_2618) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2602, input_dim2x_x1_2618, tmp_var);
      add65_2628 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2697_inst
    process(indvar_2605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2605, type_cast_2696_wire_constant, tmp_var);
      indvarx_xnext_2698 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2705_inst
    process(input_dim1x_x1x_xph_2540) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2540, type_cast_2704_wire_constant, tmp_var);
      inc_2706 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2716_inst
    process(input_dim0x_x2x_xph_2546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2546, type_cast_2715_wire_constant, tmp_var);
      inc95_2717 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2679_inst
    process(conv77_2674) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv77_2674, type_cast_2678_wire_constant, tmp_var);
      add78_2680 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2710_inst
    process(inc_2706, tmp3_2422) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2706, tmp3_2422, tmp_var);
      cmp91_2711 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2739_inst
    process(input_dim0x_x0_2735, tmp_2404) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim0x_x0_2735, tmp_2404, tmp_var);
      cmp104_2740 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2409_inst
    process(tmp_2404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2404, type_cast_2408_wire_constant, tmp_var);
      div_2410 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2427_inst
    process(tmp3_2422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2422, type_cast_2426_wire_constant, tmp_var);
      div5_2428 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2722_inst
    process(tmp3_2422) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2422, type_cast_2721_wire_constant, tmp_var);
      div98_2723 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2637_inst
    process(conv68_2632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv68_2632, type_cast_2636_wire_constant, tmp_var);
      shr118_2638 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2658_inst
    process(conv71_2653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv71_2653, type_cast_2657_wire_constant, tmp_var);
      shr72120_2659 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2556_inst
    process(tmp3_2422, input_dim0x_x2x_xph_2546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_2422, input_dim0x_x2x_xph_2546, tmp_var);
      tmp134_2557 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2566_inst
    process(tmp16_2440, tmp135_2562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2440, tmp135_2562, tmp_var);
      tmp136_2567 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2571_inst
    process(tmp41_2475, input_dim1x_x1x_xph_2540) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp41_2475, input_dim1x_x1x_xph_2540, tmp_var);
      tmp6_2572 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2581_inst
    process(tmp29_2450, input_dim0x_x2x_xph_2546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp29_2450, input_dim0x_x2x_xph_2546, tmp_var);
      tmp10_2582 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2591_inst
    process(tmp58_2511, tmp11_2587) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp58_2511, tmp11_2587, tmp_var);
      tmp12_2592 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2601_inst
    process(tmp54_2499, tmp13_2597) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_2499, tmp13_2597, tmp_var);
      tmp14_2602 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2617_inst
    process(indvar_2605) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2605, type_cast_2616_wire_constant, tmp_var);
      input_dim2x_x1_2618 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2525_inst
    process(tmp4_2521, tmp35_2465) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2521, tmp35_2465, tmp_var);
      tmp5_2526 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2536_inst
    process(tmp8_2532, tmp35_2465) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp8_2532, tmp35_2465, tmp_var);
      tmp9_2537 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2684_inst
    process(add78_2680, conv80_2515) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add78_2680, conv80_2515, tmp_var);
      cmp_2685 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2643_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr118_2642_scaled;
      array_obj_ref_2643_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2643_index_offset_req_0;
      array_obj_ref_2643_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2643_index_offset_req_1;
      array_obj_ref_2643_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2664_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr72120_2663_scaled;
      array_obj_ref_2664_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2664_index_offset_req_0;
      array_obj_ref_2664_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2664_index_offset_req_1;
      array_obj_ref_2664_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : LOAD_padding_2464_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2464_load_0_req_0;
      LOAD_padding_2464_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2464_load_0_req_1;
      LOAD_padding_2464_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2464_word_address_0;
      LOAD_padding_2464_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2421_load_0 ptr_deref_2439_load_0 ptr_deref_2403_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2421_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2439_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2403_load_0_req_0;
      ptr_deref_2421_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2439_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2403_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2421_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2439_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2403_load_0_req_1;
      ptr_deref_2421_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2439_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2403_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2421_word_address_0 & ptr_deref_2439_word_address_0 & ptr_deref_2403_word_address_0;
      ptr_deref_2421_data_0 <= data_out(47 downto 32);
      ptr_deref_2439_data_0 <= data_out(31 downto 16);
      ptr_deref_2403_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2449_load_0 ptr_deref_2474_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2449_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2474_load_0_req_0;
      ptr_deref_2449_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2474_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2449_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2474_load_0_req_1;
      ptr_deref_2449_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2474_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2449_word_address_0 & ptr_deref_2474_word_address_0;
      ptr_deref_2449_data_0 <= data_out(31 downto 16);
      ptr_deref_2474_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2486_load_0 ptr_deref_2461_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2486_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2461_load_0_req_0;
      ptr_deref_2486_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2461_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2486_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2461_load_0_req_1;
      ptr_deref_2486_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2461_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2486_word_address_0 & ptr_deref_2461_word_address_0;
      ptr_deref_2486_data_0 <= data_out(31 downto 16);
      ptr_deref_2461_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2510_load_0 ptr_deref_2498_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2510_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2498_load_0_req_0;
      ptr_deref_2510_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2498_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2510_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2498_load_0_req_1;
      ptr_deref_2510_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2498_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2510_word_address_0 & ptr_deref_2498_word_address_0;
      ptr_deref_2510_data_0 <= data_out(31 downto 16);
      ptr_deref_2498_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2648_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2648_load_0_req_0;
      ptr_deref_2648_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2648_load_0_req_1;
      ptr_deref_2648_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2648_word_address_0;
      ptr_deref_2648_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2668_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2668_store_0_req_0;
      ptr_deref_2668_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2668_store_0_req_1;
      ptr_deref_2668_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2668_word_address_0;
      data_in <= ptr_deref_2668_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2390_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2390_inst_req_0;
      RPIPE_Block3_start_2390_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2390_inst_req_1;
      RPIPE_Block3_start_2390_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2391 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2749_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2749_inst_req_0;
      WPIPE_Block3_done_2749_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2749_inst_req_1;
      WPIPE_Block3_done_2749_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2391;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_2962_start: Boolean;
  signal sendOutput_CP_2962_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1164_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1176_inst_ack_0 : boolean;
  signal if_stmt_1211_branch_ack_1 : boolean;
  signal phi_stmt_1083_req_0 : boolean;
  signal type_cast_1164_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1182_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1176_inst_req_0 : boolean;
  signal type_cast_1154_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1182_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1176_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0 : boolean;
  signal if_stmt_1211_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1182_inst_ack_0 : boolean;
  signal ptr_deref_985_load_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1197_inst_ack_1 : boolean;
  signal ptr_deref_985_load_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1176_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_req_1 : boolean;
  signal if_stmt_1211_branch_ack_0 : boolean;
  signal type_cast_1164_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1182_inst_ack_1 : boolean;
  signal type_cast_1164_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1185_inst_ack_1 : boolean;
  signal ptr_deref_985_load_0_req_1 : boolean;
  signal type_cast_989_inst_req_1 : boolean;
  signal type_cast_989_inst_ack_1 : boolean;
  signal ptr_deref_985_load_0_ack_1 : boolean;
  signal type_cast_1154_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1179_inst_req_1 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1197_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1179_inst_ack_1 : boolean;
  signal ptr_deref_1001_load_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1197_inst_req_0 : boolean;
  signal ptr_deref_1001_load_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1185_inst_ack_0 : boolean;
  signal ptr_deref_1001_load_0_req_1 : boolean;
  signal ptr_deref_1001_load_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1197_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1185_inst_req_1 : boolean;
  signal type_cast_989_inst_ack_0 : boolean;
  signal type_cast_989_inst_req_0 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1185_inst_req_0 : boolean;
  signal ptr_deref_1017_load_0_req_0 : boolean;
  signal ptr_deref_1017_load_0_ack_0 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal ptr_deref_1017_load_0_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1194_inst_ack_1 : boolean;
  signal ptr_deref_1017_load_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1194_inst_req_1 : boolean;
  signal type_cast_1154_inst_ack_0 : boolean;
  signal type_cast_1021_inst_req_0 : boolean;
  signal type_cast_1021_inst_ack_0 : boolean;
  signal type_cast_1021_inst_req_1 : boolean;
  signal type_cast_1021_inst_ack_1 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal if_stmt_1039_branch_req_0 : boolean;
  signal if_stmt_1039_branch_ack_1 : boolean;
  signal if_stmt_1039_branch_ack_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal phi_stmt_1083_ack_0 : boolean;
  signal type_cast_1066_inst_req_0 : boolean;
  signal type_cast_1066_inst_ack_0 : boolean;
  signal type_cast_1066_inst_req_1 : boolean;
  signal type_cast_1066_inst_ack_1 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1194_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1194_inst_req_0 : boolean;
  signal type_cast_1154_inst_req_0 : boolean;
  signal array_obj_ref_1095_index_offset_req_0 : boolean;
  signal array_obj_ref_1095_index_offset_ack_0 : boolean;
  signal array_obj_ref_1095_index_offset_req_1 : boolean;
  signal phi_stmt_1083_req_1 : boolean;
  signal array_obj_ref_1095_index_offset_ack_1 : boolean;
  signal type_cast_1089_inst_ack_1 : boolean;
  signal type_cast_1089_inst_req_1 : boolean;
  signal addr_of_1096_final_reg_req_0 : boolean;
  signal addr_of_1096_final_reg_ack_0 : boolean;
  signal addr_of_1096_final_reg_req_1 : boolean;
  signal addr_of_1096_final_reg_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1179_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1179_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1191_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1191_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1191_inst_ack_0 : boolean;
  signal type_cast_1089_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1191_inst_req_0 : boolean;
  signal type_cast_1089_inst_req_0 : boolean;
  signal ptr_deref_1100_load_0_req_0 : boolean;
  signal ptr_deref_1100_load_0_ack_0 : boolean;
  signal ptr_deref_1100_load_0_req_1 : boolean;
  signal ptr_deref_1100_load_0_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal type_cast_1114_inst_req_0 : boolean;
  signal type_cast_1114_inst_ack_0 : boolean;
  signal type_cast_1114_inst_req_1 : boolean;
  signal type_cast_1114_inst_ack_1 : boolean;
  signal type_cast_1124_inst_req_0 : boolean;
  signal type_cast_1124_inst_ack_0 : boolean;
  signal type_cast_1124_inst_req_1 : boolean;
  signal type_cast_1124_inst_ack_1 : boolean;
  signal type_cast_1134_inst_req_0 : boolean;
  signal type_cast_1134_inst_ack_0 : boolean;
  signal type_cast_1134_inst_req_1 : boolean;
  signal type_cast_1134_inst_ack_1 : boolean;
  signal type_cast_1144_inst_req_0 : boolean;
  signal type_cast_1144_inst_ack_0 : boolean;
  signal type_cast_1144_inst_req_1 : boolean;
  signal type_cast_1144_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_2962_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2962_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_2962_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2962_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_2962: Block -- control-path 
    signal sendOutput_CP_2962_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    sendOutput_CP_2962_elements(0) <= sendOutput_CP_2962_start;
    sendOutput_CP_2962_symbol <= sendOutput_CP_2962_elements(72);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (92) 
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/branch_block_stmt_974__entry__
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_update_start_
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Update/cr
      -- 
    rr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_985_load_0_req_0); -- 
    cr_3036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_985_load_0_req_1); -- 
    cr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => type_cast_989_inst_req_1); -- 
    rr_3089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_1001_load_0_req_0); -- 
    cr_3100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_1001_load_0_req_1); -- 
    cr_3119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => type_cast_1005_inst_req_1); -- 
    rr_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_1017_load_0_req_0); -- 
    cr_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => ptr_deref_1017_load_0_req_1); -- 
    cr_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(0), ack => type_cast_1021_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Sample/word_access_start/word_0/$exit
      -- 
    ra_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_load_0_ack_0, ack => sendOutput_CP_2962_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/ptr_deref_985_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/ptr_deref_985_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/ptr_deref_985_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/ptr_deref_985_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_985_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Sample/rr
      -- 
    ca_3037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_load_0_ack_1, ack => sendOutput_CP_2962_elements(2)); -- 
    rr_3050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(2), ack => type_cast_989_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Sample/$exit
      -- 
    ra_3051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_989_inst_ack_0, ack => sendOutput_CP_2962_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	13 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_989_update_completed_
      -- 
    ca_3056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_989_inst_ack_1, ack => sendOutput_CP_2962_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Sample/word_access_start/word_0/ra
      -- 
    ra_3090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1001_load_0_ack_0, ack => sendOutput_CP_2962_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/ptr_deref_1001_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/ptr_deref_1001_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/ptr_deref_1001_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/ptr_deref_1001_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1001_Update/word_access_complete/word_0/ca
      -- 
    ca_3101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1001_load_0_ack_1, ack => sendOutput_CP_2962_elements(6)); -- 
    rr_3114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(6), ack => type_cast_1005_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Sample/ra
      -- 
    ra_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => sendOutput_CP_2962_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1005_Update/ca
      -- 
    ca_3120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => sendOutput_CP_2962_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Sample/word_access_start/word_0/ra
      -- 
    ra_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1017_load_0_ack_0, ack => sendOutput_CP_2962_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/ptr_deref_1017_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/ptr_deref_1017_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/ptr_deref_1017_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/ptr_deref_1017_Update/ptr_deref_1017_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Sample/rr
      -- 
    ca_3165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1017_load_0_ack_1, ack => sendOutput_CP_2962_elements(10)); -- 
    rr_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(10), ack => type_cast_1021_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Sample/ra
      -- 
    ra_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1021_inst_ack_0, ack => sendOutput_CP_2962_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/type_cast_1021_Update/ca
      -- 
    ca_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1021_inst_ack_1, ack => sendOutput_CP_2962_elements(12)); -- 
    -- CP-element group 13:  branch  join  transition  place  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	4 
    -- CP-element group 13: 	8 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (10) 
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039__entry__
      -- CP-element group 13: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038__exit__
      -- CP-element group 13: 	 branch_block_stmt_974/assign_stmt_982_to_assign_stmt_1038/$exit
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_974/R_cmp77_1040_place
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_974/if_stmt_1039_else_link/$entry
      -- 
    branch_req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(13), ack => if_stmt_1039_branch_req_0); -- 
    sendOutput_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(4) & sendOutput_CP_2962_elements(8) & sendOutput_CP_2962_elements(12);
      gj_sendOutput_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (18) 
      -- CP-element group 14: 	 branch_block_stmt_974/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_974/merge_stmt_1045_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080__entry__
      -- CP-element group 14: 	 branch_block_stmt_974/merge_stmt_1045__exit__
      -- CP-element group 14: 	 branch_block_stmt_974/merge_stmt_1045_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_974/merge_stmt_1045_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_974/merge_stmt_1045_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_974/if_stmt_1039_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_974/if_stmt_1039_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_974/entry_bbx_xnph
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/$entry
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_update_start_
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_974/entry_bbx_xnph_PhiReq/$exit
      -- 
    if_choice_transition_3197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_1, ack => sendOutput_CP_2962_elements(14)); -- 
    rr_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(14), ack => type_cast_1066_inst_req_0); -- 
    cr_3219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(14), ack => type_cast_1066_inst_req_1); -- 
    -- CP-element group 15:  transition  place  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	72 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_974/entry_forx_xend_PhiReq/$exit
      -- CP-element group 15: 	 branch_block_stmt_974/entry_forx_xend_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_974/if_stmt_1039_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_974/if_stmt_1039_else_link/else_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_974/entry_forx_xend
      -- 
    else_choice_transition_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1039_branch_ack_0, ack => sendOutput_CP_2962_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Sample/ra
      -- 
    ra_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_0, ack => sendOutput_CP_2962_elements(16)); -- 
    -- CP-element group 17:  transition  place  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	66 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080__exit__
      -- CP-element group 17: 	 branch_block_stmt_974/bbx_xnph_forx_xbody
      -- CP-element group 17: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/$entry
      -- CP-element group 17: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/$exit
      -- CP-element group 17: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_974/assign_stmt_1051_to_assign_stmt_1080/type_cast_1066_Update/ca
      -- 
    ca_3220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1066_inst_ack_1, ack => sendOutput_CP_2962_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	71 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	63 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Sample/ack
      -- 
    ack_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1095_index_offset_ack_0, ack => sendOutput_CP_2962_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	71 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (11) 
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_root_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_offset_calculated
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_base_plus_offset/$entry
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_base_plus_offset/$exit
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_request/$entry
      -- CP-element group 19: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_request/req
      -- 
    ack_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1095_index_offset_ack_1, ack => sendOutput_CP_2962_elements(19)); -- 
    req_3263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(19), ack => addr_of_1096_final_reg_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_request/$exit
      -- CP-element group 20: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_request/ack
      -- 
    ack_3264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1096_final_reg_ack_0, ack => sendOutput_CP_2962_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	71 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (24) 
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_complete/ack
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_word_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_root_address_calculated
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_address_resized
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_addr_resize/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_addr_resize/$exit
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_plus_offset/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_plus_offset/$exit
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_word_addrgen/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_word_addrgen/$exit
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_word_addrgen/root_register_req
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_word_addrgen/root_register_ack
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/word_0/$entry
      -- CP-element group 21: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/word_0/rr
      -- 
    ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1096_final_reg_ack_1, ack => sendOutput_CP_2962_elements(21)); -- 
    rr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(21), ack => ptr_deref_1100_load_0_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/$exit
      -- CP-element group 22: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Sample/word_access_start/word_0/ra
      -- 
    ra_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1100_load_0_ack_0, ack => sendOutput_CP_2962_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	71 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	26 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	34 
    -- CP-element group 23: 	36 
    -- CP-element group 23: 	38 
    -- CP-element group 23:  members (33) 
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/$exit
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/word_0/ca
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/ptr_deref_1100_Merge/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/ptr_deref_1100_Merge/$exit
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/ptr_deref_1100_Merge/merge_req
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/ptr_deref_1100_Merge/merge_ack
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_sample_start_
      -- 
    ca_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1100_load_0_ack_1, ack => sendOutput_CP_2962_elements(23)); -- 
    rr_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1124_inst_req_0); -- 
    rr_3369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1134_inst_req_0); -- 
    rr_3383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1144_inst_req_0); -- 
    rr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1104_inst_req_0); -- 
    rr_3341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1114_inst_req_0); -- 
    rr_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1154_inst_req_0); -- 
    rr_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1164_inst_req_0); -- 
    rr_3425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(23), ack => type_cast_1174_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Sample/ra
      -- 
    ra_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => sendOutput_CP_2962_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	71 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	60 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Update/ca
      -- 
    ca_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => sendOutput_CP_2962_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Sample/ra
      -- 
    ra_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1114_inst_ack_0, ack => sendOutput_CP_2962_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	71 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	57 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Update/ca
      -- 
    ca_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1114_inst_ack_1, ack => sendOutput_CP_2962_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Sample/ra
      -- 
    ra_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1124_inst_ack_0, ack => sendOutput_CP_2962_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	71 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	54 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Update/ca
      -- 
    ca_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1124_inst_ack_1, ack => sendOutput_CP_2962_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Sample/ra
      -- 
    ra_3370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_0, ack => sendOutput_CP_2962_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	71 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	51 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Update/ca
      -- 
    ca_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_1, ack => sendOutput_CP_2962_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Sample/ra
      -- 
    ra_3384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_0, ack => sendOutput_CP_2962_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	71 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	48 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Update/ca
      -- 
    ca_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1144_inst_ack_1, ack => sendOutput_CP_2962_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_sample_completed_
      -- 
    ra_3398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1154_inst_ack_0, ack => sendOutput_CP_2962_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	71 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	45 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_update_completed_
      -- 
    ca_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1154_inst_ack_1, ack => sendOutput_CP_2962_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	23 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Sample/$exit
      -- 
    ra_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_0, ack => sendOutput_CP_2962_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	71 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	42 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_update_completed_
      -- 
    ca_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_1, ack => sendOutput_CP_2962_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	23 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Sample/$exit
      -- 
    ra_3426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => sendOutput_CP_2962_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	71 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Sample/req
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_update_completed_
      -- 
    ca_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => sendOutput_CP_2962_elements(39)); -- 
    req_3439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1176_inst_req_0); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Update/req
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_update_start_
      -- CP-element group 40: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Update/$entry
      -- 
    ack_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1176_inst_ack_0, ack => sendOutput_CP_2962_elements(40)); -- 
    req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1176_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1176_update_completed_
      -- 
    ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1176_inst_ack_1, ack => sendOutput_CP_2962_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	37 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Sample/$entry
      -- 
    req_3453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1179_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(41) & sendOutput_CP_2962_elements(37);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Update/req
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_update_start_
      -- 
    ack_3454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1179_inst_ack_0, ack => sendOutput_CP_2962_elements(43)); -- 
    req_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1179_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1179_update_completed_
      -- 
    ack_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1179_inst_ack_1, ack => sendOutput_CP_2962_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	35 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Sample/req
      -- CP-element group 45: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_sample_start_
      -- 
    req_3467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1182_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(44) & sendOutput_CP_2962_elements(35);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Update/req
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_update_start_
      -- 
    ack_3468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1182_inst_ack_0, ack => sendOutput_CP_2962_elements(46)); -- 
    req_3472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1182_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1182_update_completed_
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1182_inst_ack_1, ack => sendOutput_CP_2962_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	33 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Sample/req
      -- CP-element group 48: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_sample_start_
      -- 
    req_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1185_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(33) & sendOutput_CP_2962_elements(47);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Update/req
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_update_start_
      -- CP-element group 49: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_sample_completed_
      -- 
    ack_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1185_inst_ack_0, ack => sendOutput_CP_2962_elements(49)); -- 
    req_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1185_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1185_update_completed_
      -- 
    ack_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1185_inst_ack_1, ack => sendOutput_CP_2962_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	31 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Sample/$entry
      -- 
    req_3495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1188_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(31) & sendOutput_CP_2962_elements(50);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_update_start_
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Update/req
      -- CP-element group 52: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_sample_completed_
      -- 
    ack_3496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0, ack => sendOutput_CP_2962_elements(52)); -- 
    req_3500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1188_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1188_Update/ack
      -- 
    ack_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1, ack => sendOutput_CP_2962_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	29 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_sample_start_
      -- 
    req_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1191_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(29) & sendOutput_CP_2962_elements(53);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Update/req
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_update_start_
      -- CP-element group 55: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_sample_completed_
      -- 
    ack_3510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1191_inst_ack_0, ack => sendOutput_CP_2962_elements(55)); -- 
    req_3514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1191_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1191_update_completed_
      -- 
    ack_3515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1191_inst_ack_1, ack => sendOutput_CP_2962_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	27 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Sample/req
      -- CP-element group 57: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_sample_start_
      -- 
    req_3523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(57), ack => WPIPE_ConvTranspose_output_pipe_1194_inst_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(27) & sendOutput_CP_2962_elements(56);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Update/req
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_update_start_
      -- CP-element group 58: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_sample_completed_
      -- 
    ack_3524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1194_inst_ack_0, ack => sendOutput_CP_2962_elements(58)); -- 
    req_3528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(58), ack => WPIPE_ConvTranspose_output_pipe_1194_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1194_update_completed_
      -- 
    ack_3529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1194_inst_ack_1, ack => sendOutput_CP_2962_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	25 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_sample_start_
      -- 
    req_3537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(60), ack => WPIPE_ConvTranspose_output_pipe_1197_inst_req_0); -- 
    sendOutput_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(25) & sendOutput_CP_2962_elements(59);
      gj_sendOutput_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Update/req
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_update_start_
      -- CP-element group 61: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_sample_completed_
      -- 
    ack_3538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1197_inst_ack_0, ack => sendOutput_CP_2962_elements(61)); -- 
    req_3542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(61), ack => WPIPE_ConvTranspose_output_pipe_1197_inst_req_1); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/WPIPE_ConvTranspose_output_pipe_1197_update_completed_
      -- 
    ack_3543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1197_inst_ack_1, ack => sendOutput_CP_2962_elements(62)); -- 
    -- CP-element group 63:  branch  join  transition  place  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	18 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (10) 
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_if_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_eval_test/branch_req
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_eval_test/$entry
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_else_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210__exit__
      -- CP-element group 63: 	 branch_block_stmt_974/R_exitcond1_1212_place
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211__entry__
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_eval_test/$exit
      -- CP-element group 63: 	 branch_block_stmt_974/if_stmt_1211_dead_link/$entry
      -- CP-element group 63: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/$exit
      -- 
    branch_req_3551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(63), ack => if_stmt_1211_branch_req_0); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(18) & sendOutput_CP_2962_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	72 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_974/merge_stmt_1217_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_974/if_stmt_1211_if_link/if_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 64: 	 branch_block_stmt_974/if_stmt_1211_if_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_974/merge_stmt_1217__exit__
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xendx_xloopexit_forx_xend
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_974/merge_stmt_1217_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_974/merge_stmt_1217_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_974/merge_stmt_1217_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_974/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_3556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1211_branch_ack_1, ack => sendOutput_CP_2962_elements(64)); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (12) 
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/if_stmt_1211_else_link/else_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_974/if_stmt_1211_else_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Update/cr
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1211_branch_ack_0, ack => sendOutput_CP_2962_elements(65)); -- 
    cr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(65), ack => type_cast_1089_inst_req_1); -- 
    rr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(65), ack => type_cast_1089_inst_req_0); -- 
    -- CP-element group 66:  transition  output  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	17 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	70 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_req
      -- CP-element group 66: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1087_konst_delay_trans
      -- CP-element group 66: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1083/$exit
      -- CP-element group 66: 	 branch_block_stmt_974/bbx_xnph_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_1083_req_3585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1083_req_3585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(66), ack => phi_stmt_1083_req_0); -- 
    -- Element group sendOutput_CP_2962_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => sendOutput_CP_2962_elements(17), ack => sendOutput_CP_2962_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Sample/$exit
      -- 
    ra_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_0, ack => sendOutput_CP_2962_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Update/ca
      -- CP-element group 68: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/Update/$exit
      -- 
    ca_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1089_inst_ack_1, ack => sendOutput_CP_2962_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/$exit
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/$exit
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_sources/type_cast_1089/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_974/forx_xbody_forx_xbody_PhiReq/phi_stmt_1083/phi_stmt_1083_req
      -- 
    phi_stmt_1083_req_3611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1083_req_3611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(69), ack => phi_stmt_1083_req_1); -- 
    sendOutput_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2962_elements(67) & sendOutput_CP_2962_elements(68);
      gj_sendOutput_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2962_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  merge  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	66 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_974/merge_stmt_1082_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_974/merge_stmt_1082_PhiAck/$entry
      -- 
    sendOutput_CP_2962_elements(70) <= OrReduce(sendOutput_CP_2962_elements(66) & sendOutput_CP_2962_elements(69));
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	27 
    -- CP-element group 71: 	29 
    -- CP-element group 71: 	31 
    -- CP-element group 71: 	39 
    -- CP-element group 71: 	25 
    -- CP-element group 71: 	33 
    -- CP-element group 71: 	35 
    -- CP-element group 71: 	37 
    -- CP-element group 71: 	23 
    -- CP-element group 71: 	21 
    -- CP-element group 71: 	18 
    -- CP-element group 71: 	19 
    -- CP-element group 71:  members (53) 
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1164_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210__entry__
      -- CP-element group 71: 	 branch_block_stmt_974/merge_stmt_1082__exit__
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/merge_stmt_1082_PhiAck/phi_stmt_1083_ack
      -- CP-element group 71: 	 branch_block_stmt_974/merge_stmt_1082_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_resized_1
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_scaled_1
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_computed_1
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1174_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_resize_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_resize_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_resize_1/index_resize_req
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_resize_1/index_resize_ack
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_scale_1/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_scale_1/$exit
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_scale_1/scale_rename_req
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_index_scale_1/scale_rename_ack
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/array_obj_ref_1095_final_index_sum_regn_Update/req
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_complete/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/addr_of_1096_complete/req
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/word_0/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/ptr_deref_1100_Update/word_access_complete/word_0/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1104_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1114_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1124_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1134_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_update_start_
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1144_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_974/assign_stmt_1097_to_assign_stmt_1210/type_cast_1154_update_start_
      -- 
    phi_stmt_1083_ack_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1083_ack_0, ack => sendOutput_CP_2962_elements(71)); -- 
    cr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1164_inst_req_1); -- 
    cr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1154_inst_req_1); -- 
    cr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1174_inst_req_1); -- 
    req_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => array_obj_ref_1095_index_offset_req_0); -- 
    req_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => array_obj_ref_1095_index_offset_req_1); -- 
    req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => addr_of_1096_final_reg_req_1); -- 
    cr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => ptr_deref_1100_load_0_req_1); -- 
    cr_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1104_inst_req_1); -- 
    cr_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1114_inst_req_1); -- 
    cr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1124_inst_req_1); -- 
    cr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1134_inst_req_1); -- 
    cr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2962_elements(71), ack => type_cast_1144_inst_req_1); -- 
    -- CP-element group 72:  merge  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	15 
    -- CP-element group 72: 	64 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1219_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_974/branch_block_stmt_974__exit__
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1221_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1221__exit__
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1219__exit__
      -- CP-element group 72: 	 branch_block_stmt_974/return__
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1221_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_974/$exit
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1219_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1221_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1221_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1219_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_974/merge_stmt_1219_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_974/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_974/return___PhiReq/$entry
      -- 
    sendOutput_CP_2962_elements(72) <= OrReduce(sendOutput_CP_2962_elements(15) & sendOutput_CP_2962_elements(64));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1094_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1094_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1095_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1097 : std_logic_vector(31 downto 0);
    signal cmp77_1038 : std_logic_vector(0 downto 0);
    signal conv15_1105 : std_logic_vector(7 downto 0);
    signal conv21_1115 : std_logic_vector(7 downto 0);
    signal conv27_1125 : std_logic_vector(7 downto 0);
    signal conv2_1006 : std_logic_vector(31 downto 0);
    signal conv33_1135 : std_logic_vector(7 downto 0);
    signal conv39_1145 : std_logic_vector(7 downto 0);
    signal conv45_1155 : std_logic_vector(7 downto 0);
    signal conv4_1022 : std_logic_vector(31 downto 0);
    signal conv51_1165 : std_logic_vector(7 downto 0);
    signal conv57_1175 : std_logic_vector(7 downto 0);
    signal conv_990 : std_logic_vector(31 downto 0);
    signal exitcond1_1210 : std_logic_vector(0 downto 0);
    signal iNsTr_0_982 : std_logic_vector(31 downto 0);
    signal iNsTr_1_998 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1014 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1067 : std_logic_vector(63 downto 0);
    signal indvar_1083 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1205 : std_logic_vector(63 downto 0);
    signal mul5_1032 : std_logic_vector(31 downto 0);
    signal mul_1027 : std_logic_vector(31 downto 0);
    signal ptr_deref_1001_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1001_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1001_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1001_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1001_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1017_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1017_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1017_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1017_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1017_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1100_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1100_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1100_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1100_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1100_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_985_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_985_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_985_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_985_word_offset_0 : std_logic_vector(6 downto 0);
    signal shr18_1111 : std_logic_vector(63 downto 0);
    signal shr24_1121 : std_logic_vector(63 downto 0);
    signal shr30_1131 : std_logic_vector(63 downto 0);
    signal shr36_1141 : std_logic_vector(63 downto 0);
    signal shr42_1151 : std_logic_vector(63 downto 0);
    signal shr48_1161 : std_logic_vector(63 downto 0);
    signal shr54_1171 : std_logic_vector(63 downto 0);
    signal tmp12_1101 : std_logic_vector(63 downto 0);
    signal tmp1_1002 : std_logic_vector(15 downto 0);
    signal tmp3_1018 : std_logic_vector(15 downto 0);
    signal tmp84_1051 : std_logic_vector(31 downto 0);
    signal tmp84x_xop_1063 : std_logic_vector(31 downto 0);
    signal tmp85_1057 : std_logic_vector(0 downto 0);
    signal tmp88_1080 : std_logic_vector(63 downto 0);
    signal tmp_986 : std_logic_vector(15 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1071_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1087_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1089_wire : std_logic_vector(63 downto 0);
    signal type_cast_1109_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1119_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1129_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1139_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1159_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1169_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1073 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1095_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1095_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1095_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1095_resized_base_address <= "00000000000000";
    iNsTr_0_982 <= "00000000000000000000000000000011";
    iNsTr_1_998 <= "00000000000000000000000000000100";
    iNsTr_2_1014 <= "00000000000000000000000000000101";
    ptr_deref_1001_word_offset_0 <= "0000000";
    ptr_deref_1017_word_offset_0 <= "0000000";
    ptr_deref_1100_word_offset_0 <= "00000000000000";
    ptr_deref_985_word_offset_0 <= "0000000";
    type_cast_1036_wire_constant <= "00000000000000000000000000000011";
    type_cast_1049_wire_constant <= "00000000000000000000000000000010";
    type_cast_1055_wire_constant <= "00000000000000000000000000000001";
    type_cast_1061_wire_constant <= "11111111111111111111111111111111";
    type_cast_1071_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1087_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1109_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1119_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1129_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1139_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1149_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1159_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1169_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1083: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1087_wire_constant & type_cast_1089_wire;
      req <= phi_stmt_1083_req_0 & phi_stmt_1083_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1083",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1083_ack_0,
          idata => idata,
          odata => indvar_1083,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1083
    -- flow-through select operator MUX_1079_inst
    tmp88_1080 <= xx_xop_1073 when (tmp85_1057(0) /=  '0') else type_cast_1078_wire_constant;
    addr_of_1096_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1096_final_reg_req_0;
      addr_of_1096_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1096_final_reg_req_1;
      addr_of_1096_final_reg_ack_1<= rack(0);
      addr_of_1096_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1096_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1095_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1097,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1002,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_1006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1021_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1021_inst_req_0;
      type_cast_1021_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1021_inst_req_1;
      type_cast_1021_inst_ack_1<= rack(0);
      type_cast_1021_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1021_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_1022,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1066_inst_req_0;
      type_cast_1066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1066_inst_req_1;
      type_cast_1066_inst_ack_1<= rack(0);
      type_cast_1066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp84x_xop_1063,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1089_inst_req_0;
      type_cast_1089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1089_inst_req_1;
      type_cast_1089_inst_ack_1<= rack(0);
      type_cast_1089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1089_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1114_inst_req_0;
      type_cast_1114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1114_inst_req_1;
      type_cast_1114_inst_ack_1<= rack(0);
      type_cast_1114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr18_1111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_1115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1124_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1124_inst_req_0;
      type_cast_1124_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1124_inst_req_1;
      type_cast_1124_inst_ack_1<= rack(0);
      type_cast_1124_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1124_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr24_1121,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1125,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1134_inst_req_0;
      type_cast_1134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1134_inst_req_1;
      type_cast_1134_inst_ack_1<= rack(0);
      type_cast_1134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr30_1131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1144_inst_req_0;
      type_cast_1144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1144_inst_req_1;
      type_cast_1144_inst_ack_1<= rack(0);
      type_cast_1144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr36_1141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1154_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1154_inst_req_0;
      type_cast_1154_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1154_inst_req_1;
      type_cast_1154_inst_ack_1<= rack(0);
      type_cast_1154_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1154_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr42_1151,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_1155,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1164_inst_req_0;
      type_cast_1164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1164_inst_req_1;
      type_cast_1164_inst_ack_1<= rack(0);
      type_cast_1164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr48_1161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_1165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr54_1171,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_989_inst_req_0;
      type_cast_989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_989_inst_req_1;
      type_cast_989_inst_ack_1<= rack(0);
      type_cast_989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_989_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_986,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_990,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1095_index_1_rename
    process(R_indvar_1094_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1094_resized;
      ov(13 downto 0) := iv;
      R_indvar_1094_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1095_index_1_resize
    process(indvar_1083) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1083;
      ov := iv(13 downto 0);
      R_indvar_1094_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1095_root_address_inst
    process(array_obj_ref_1095_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1095_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1095_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1001_addr_0
    process(ptr_deref_1001_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1001_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1001_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1001_base_resize
    process(iNsTr_1_998) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_998;
      ov := iv(6 downto 0);
      ptr_deref_1001_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1001_gather_scatter
    process(ptr_deref_1001_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1001_data_0;
      ov(15 downto 0) := iv;
      tmp1_1002 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1001_root_address_inst
    process(ptr_deref_1001_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1001_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1001_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1017_addr_0
    process(ptr_deref_1017_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1017_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1017_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1017_base_resize
    process(iNsTr_2_1014) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1014;
      ov := iv(6 downto 0);
      ptr_deref_1017_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1017_gather_scatter
    process(ptr_deref_1017_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1017_data_0;
      ov(15 downto 0) := iv;
      tmp3_1018 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1017_root_address_inst
    process(ptr_deref_1017_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1017_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1017_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1100_addr_0
    process(ptr_deref_1100_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1100_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1100_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1100_base_resize
    process(arrayidx_1097) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1097;
      ov := iv(13 downto 0);
      ptr_deref_1100_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1100_gather_scatter
    process(ptr_deref_1100_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1100_data_0;
      ov(63 downto 0) := iv;
      tmp12_1101 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1100_root_address_inst
    process(ptr_deref_1100_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1100_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1100_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_985_addr_0
    process(ptr_deref_985_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_985_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_985_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_985_base_resize
    process(iNsTr_0_982) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_982;
      ov := iv(6 downto 0);
      ptr_deref_985_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_985_gather_scatter
    process(ptr_deref_985_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_985_data_0;
      ov(15 downto 0) := iv;
      tmp_986 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_985_root_address_inst
    process(ptr_deref_985_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_985_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_985_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1039_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1038;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1039_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1039_branch_req_0,
          ack0 => if_stmt_1039_branch_ack_0,
          ack1 => if_stmt_1039_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1211_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1210;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1211_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1211_branch_req_0,
          ack0 => if_stmt_1211_branch_ack_0,
          ack1 => if_stmt_1211_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1062_inst
    process(tmp84_1051) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp84_1051, type_cast_1061_wire_constant, tmp_var);
      tmp84x_xop_1063 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1072_inst
    process(iNsTr_4_1067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1067, type_cast_1071_wire_constant, tmp_var);
      xx_xop_1073 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1204_inst
    process(indvar_1083) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1083, type_cast_1203_wire_constant, tmp_var);
      indvarx_xnext_1205 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1209_inst
    process(indvarx_xnext_1205, tmp88_1080) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1205, tmp88_1080, tmp_var);
      exitcond1_1210 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1050_inst
    process(mul5_1032) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul5_1032, type_cast_1049_wire_constant, tmp_var);
      tmp84_1051 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1110_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1109_wire_constant, tmp_var);
      shr18_1111 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1120_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1119_wire_constant, tmp_var);
      shr24_1121 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1130_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1129_wire_constant, tmp_var);
      shr30_1131 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1140_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1139_wire_constant, tmp_var);
      shr36_1141 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1150_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1149_wire_constant, tmp_var);
      shr42_1151 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1160_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1159_wire_constant, tmp_var);
      shr48_1161 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1170_inst
    process(tmp12_1101) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp12_1101, type_cast_1169_wire_constant, tmp_var);
      shr54_1171 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1026_inst
    process(conv2_1006, conv_990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv2_1006, conv_990, tmp_var);
      mul_1027 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1031_inst
    process(mul_1027, conv4_1022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1027, conv4_1022, tmp_var);
      mul5_1032 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1037_inst
    process(mul5_1032) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul5_1032, type_cast_1036_wire_constant, tmp_var);
      cmp77_1038 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1056_inst
    process(tmp84_1051) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp84_1051, type_cast_1055_wire_constant, tmp_var);
      tmp85_1057 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1095_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1094_scaled;
      array_obj_ref_1095_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1095_index_offset_req_0;
      array_obj_ref_1095_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1095_index_offset_req_1;
      array_obj_ref_1095_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1001_load_0 ptr_deref_985_load_0 ptr_deref_1017_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1001_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_985_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1017_load_0_req_0;
      ptr_deref_1001_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_985_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1017_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1001_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_985_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1017_load_0_req_1;
      ptr_deref_1001_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_985_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1017_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1001_word_address_0 & ptr_deref_985_word_address_0 & ptr_deref_1017_word_address_0;
      ptr_deref_1001_data_0 <= data_out(47 downto 32);
      ptr_deref_985_data_0 <= data_out(31 downto 16);
      ptr_deref_1017_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1100_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1100_load_0_req_0;
      ptr_deref_1100_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1100_load_0_req_1;
      ptr_deref_1100_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1100_word_address_0;
      ptr_deref_1100_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(13 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(63 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1176_inst WPIPE_ConvTranspose_output_pipe_1179_inst WPIPE_ConvTranspose_output_pipe_1185_inst WPIPE_ConvTranspose_output_pipe_1182_inst WPIPE_ConvTranspose_output_pipe_1188_inst WPIPE_ConvTranspose_output_pipe_1191_inst WPIPE_ConvTranspose_output_pipe_1194_inst WPIPE_ConvTranspose_output_pipe_1197_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1176_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1179_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1185_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1182_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1188_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1191_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1194_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1197_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1176_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1179_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1185_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1182_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1188_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1191_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1194_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1197_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1176_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1179_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1185_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1182_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1188_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1191_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1194_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1197_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1176_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1179_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1185_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1182_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1188_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1191_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1194_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1197_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv57_1175 & conv51_1165 & conv39_1145 & conv45_1155 & conv33_1135 & conv27_1125 & conv21_1115 & conv15_1105;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_934_inst_req_1 : boolean;
  signal ptr_deref_468_load_0_ack_1 : boolean;
  signal type_cast_192_inst_ack_1 : boolean;
  signal type_cast_862_inst_ack_1 : boolean;
  signal type_cast_488_inst_req_1 : boolean;
  signal type_cast_488_inst_ack_1 : boolean;
  signal type_cast_192_inst_req_1 : boolean;
  signal phi_stmt_157_req_1 : boolean;
  signal type_cast_488_inst_req_0 : boolean;
  signal type_cast_488_inst_ack_0 : boolean;
  signal type_cast_162_inst_ack_1 : boolean;
  signal type_cast_162_inst_req_1 : boolean;
  signal ptr_deref_381_store_0_ack_0 : boolean;
  signal type_cast_398_inst_ack_1 : boolean;
  signal ptr_deref_381_store_0_req_0 : boolean;
  signal type_cast_398_inst_req_1 : boolean;
  signal type_cast_398_inst_ack_0 : boolean;
  signal type_cast_398_inst_req_0 : boolean;
  signal ptr_deref_468_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_160_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal ptr_deref_394_load_0_ack_1 : boolean;
  signal ptr_deref_394_load_0_req_1 : boolean;
  signal ptr_deref_122_load_0_req_0 : boolean;
  signal ptr_deref_122_load_0_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal ptr_deref_47_store_0_req_0 : boolean;
  signal ptr_deref_47_store_0_ack_0 : boolean;
  signal ptr_deref_47_store_0_req_1 : boolean;
  signal ptr_deref_47_store_0_ack_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_1 : boolean;
  signal ptr_deref_426_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal type_cast_62_inst_req_0 : boolean;
  signal ptr_deref_426_load_0_req_0 : boolean;
  signal type_cast_62_inst_ack_0 : boolean;
  signal type_cast_62_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_1 : boolean;
  signal type_cast_62_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_ack_1 : boolean;
  signal if_stmt_64_branch_req_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal if_stmt_64_branch_ack_1 : boolean;
  signal if_stmt_64_branch_ack_0 : boolean;
  signal type_cast_414_inst_ack_1 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal ptr_deref_484_load_0_ack_1 : boolean;
  signal type_cast_472_inst_ack_1 : boolean;
  signal type_cast_414_inst_req_1 : boolean;
  signal array_obj_ref_101_index_offset_req_0 : boolean;
  signal array_obj_ref_101_index_offset_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_1 : boolean;
  signal type_cast_160_inst_ack_1 : boolean;
  signal array_obj_ref_101_index_offset_ack_1 : boolean;
  signal ptr_deref_468_load_0_ack_0 : boolean;
  signal addr_of_102_final_reg_req_0 : boolean;
  signal addr_of_102_final_reg_ack_0 : boolean;
  signal addr_of_102_final_reg_req_1 : boolean;
  signal addr_of_102_final_reg_ack_1 : boolean;
  signal ptr_deref_484_load_0_req_1 : boolean;
  signal type_cast_430_inst_ack_1 : boolean;
  signal ptr_deref_468_load_0_req_0 : boolean;
  signal type_cast_472_inst_req_1 : boolean;
  signal ptr_deref_105_store_0_req_0 : boolean;
  signal ptr_deref_410_load_0_ack_1 : boolean;
  signal ptr_deref_105_store_0_ack_0 : boolean;
  signal ptr_deref_105_store_0_req_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal ptr_deref_105_store_0_ack_1 : boolean;
  signal type_cast_430_inst_req_1 : boolean;
  signal type_cast_430_inst_ack_0 : boolean;
  signal type_cast_430_inst_req_0 : boolean;
  signal ptr_deref_410_load_0_req_1 : boolean;
  signal ptr_deref_381_store_0_ack_1 : boolean;
  signal ptr_deref_381_store_0_req_1 : boolean;
  signal addr_of_287_final_reg_req_0 : boolean;
  signal addr_of_287_final_reg_ack_0 : boolean;
  signal addr_of_287_final_reg_req_1 : boolean;
  signal addr_of_287_final_reg_ack_1 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal ptr_deref_122_load_0_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal ptr_deref_122_load_0_ack_1 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_414_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_ack_1 : boolean;
  signal type_cast_160_inst_ack_0 : boolean;
  signal type_cast_141_inst_req_0 : boolean;
  signal type_cast_141_inst_ack_0 : boolean;
  signal type_cast_141_inst_req_1 : boolean;
  signal type_cast_141_inst_ack_1 : boolean;
  signal phi_stmt_157_ack_0 : boolean;
  signal phi_stmt_73_req_0 : boolean;
  signal if_stmt_143_branch_req_0 : boolean;
  signal if_stmt_143_branch_ack_1 : boolean;
  signal type_cast_414_inst_req_0 : boolean;
  signal if_stmt_143_branch_ack_0 : boolean;
  signal type_cast_934_inst_ack_1 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal ptr_deref_171_store_0_req_0 : boolean;
  signal ptr_deref_171_store_0_ack_0 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal ptr_deref_171_store_0_req_1 : boolean;
  signal ptr_deref_171_store_0_ack_1 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal ptr_deref_452_load_0_ack_1 : boolean;
  signal if_stmt_180_branch_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal ptr_deref_410_load_0_ack_0 : boolean;
  signal if_stmt_180_branch_ack_1 : boolean;
  signal if_stmt_180_branch_ack_0 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal ptr_deref_452_load_0_req_1 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_req_0 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_ack_0 : boolean;
  signal type_cast_472_inst_ack_0 : boolean;
  signal ptr_deref_410_load_0_req_0 : boolean;
  signal type_cast_472_inst_req_0 : boolean;
  signal array_obj_ref_211_index_offset_req_0 : boolean;
  signal array_obj_ref_211_index_offset_ack_0 : boolean;
  signal array_obj_ref_211_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 : boolean;
  signal array_obj_ref_211_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_876_inst_req_0 : boolean;
  signal addr_of_212_final_reg_req_0 : boolean;
  signal addr_of_212_final_reg_ack_0 : boolean;
  signal addr_of_212_final_reg_req_1 : boolean;
  signal addr_of_212_final_reg_ack_1 : boolean;
  signal ptr_deref_484_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_req_0 : boolean;
  signal phi_stmt_157_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_ack_1 : boolean;
  signal type_cast_160_inst_req_0 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal ptr_deref_484_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_930_inst_req_1 : boolean;
  signal ptr_deref_394_load_0_ack_0 : boolean;
  signal phi_stmt_189_req_0 : boolean;
  signal ptr_deref_394_load_0_req_0 : boolean;
  signal ptr_deref_222_store_0_req_0 : boolean;
  signal ptr_deref_222_store_0_ack_0 : boolean;
  signal ptr_deref_222_store_0_req_1 : boolean;
  signal ptr_deref_222_store_0_ack_1 : boolean;
  signal ptr_deref_239_load_0_req_0 : boolean;
  signal ptr_deref_239_load_0_ack_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal ptr_deref_239_load_0_req_1 : boolean;
  signal ptr_deref_239_load_0_ack_1 : boolean;
  signal type_cast_243_inst_req_0 : boolean;
  signal type_cast_243_inst_ack_0 : boolean;
  signal type_cast_243_inst_req_1 : boolean;
  signal type_cast_243_inst_ack_1 : boolean;
  signal ptr_deref_452_load_0_ack_0 : boolean;
  signal if_stmt_252_branch_req_0 : boolean;
  signal if_stmt_252_branch_ack_1 : boolean;
  signal if_stmt_252_branch_ack_0 : boolean;
  signal ptr_deref_452_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 : boolean;
  signal ptr_deref_426_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal ptr_deref_426_load_0_req_1 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal type_cast_898_inst_req_0 : boolean;
  signal ptr_deref_290_store_0_req_0 : boolean;
  signal ptr_deref_290_store_0_ack_0 : boolean;
  signal ptr_deref_290_store_0_req_1 : boolean;
  signal ptr_deref_290_store_0_ack_1 : boolean;
  signal type_cast_898_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 : boolean;
  signal type_cast_298_inst_req_0 : boolean;
  signal type_cast_298_inst_ack_0 : boolean;
  signal type_cast_298_inst_req_1 : boolean;
  signal type_cast_298_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal phi_stmt_80_req_1 : boolean;
  signal if_stmt_312_branch_req_0 : boolean;
  signal if_stmt_312_branch_ack_1 : boolean;
  signal if_stmt_312_branch_ack_0 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal STORE_padding_324_store_0_req_0 : boolean;
  signal STORE_padding_324_store_0_ack_0 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal STORE_padding_324_store_0_req_1 : boolean;
  signal STORE_padding_324_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 : boolean;
  signal type_cast_880_inst_req_1 : boolean;
  signal type_cast_332_inst_req_0 : boolean;
  signal type_cast_332_inst_ack_0 : boolean;
  signal type_cast_332_inst_req_1 : boolean;
  signal type_cast_332_inst_ack_1 : boolean;
  signal type_cast_880_inst_ack_1 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_934_inst_req_0 : boolean;
  signal type_cast_934_inst_ack_0 : boolean;
  signal ptr_deref_343_store_0_req_0 : boolean;
  signal ptr_deref_343_store_0_ack_0 : boolean;
  signal ptr_deref_343_store_0_req_1 : boolean;
  signal ptr_deref_343_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 : boolean;
  signal type_cast_351_inst_req_0 : boolean;
  signal type_cast_351_inst_ack_0 : boolean;
  signal type_cast_351_inst_req_1 : boolean;
  signal type_cast_351_inst_ack_1 : boolean;
  signal ptr_deref_362_store_0_req_0 : boolean;
  signal ptr_deref_362_store_0_ack_0 : boolean;
  signal ptr_deref_362_store_0_req_1 : boolean;
  signal ptr_deref_362_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 : boolean;
  signal ptr_deref_500_load_0_req_0 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal ptr_deref_500_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_894_inst_req_0 : boolean;
  signal ptr_deref_500_load_0_req_1 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal ptr_deref_500_load_0_ack_1 : boolean;
  signal type_cast_862_inst_req_1 : boolean;
  signal type_cast_504_inst_req_0 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal phi_stmt_73_req_1 : boolean;
  signal type_cast_504_inst_req_1 : boolean;
  signal type_cast_504_inst_ack_1 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal type_cast_192_inst_ack_0 : boolean;
  signal type_cast_192_inst_req_0 : boolean;
  signal if_stmt_527_branch_req_0 : boolean;
  signal if_stmt_527_branch_ack_1 : boolean;
  signal if_stmt_527_branch_ack_0 : boolean;
  signal type_cast_162_inst_ack_0 : boolean;
  signal if_stmt_542_branch_req_0 : boolean;
  signal if_stmt_542_branch_ack_1 : boolean;
  signal if_stmt_542_branch_ack_0 : boolean;
  signal phi_stmt_80_req_0 : boolean;
  signal type_cast_569_inst_req_0 : boolean;
  signal type_cast_569_inst_ack_0 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal type_cast_569_inst_req_1 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal type_cast_569_inst_ack_1 : boolean;
  signal if_stmt_956_branch_ack_0 : boolean;
  signal phi_stmt_189_ack_0 : boolean;
  signal array_obj_ref_598_index_offset_req_0 : boolean;
  signal array_obj_ref_598_index_offset_ack_0 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal array_obj_ref_598_index_offset_req_1 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal array_obj_ref_598_index_offset_ack_1 : boolean;
  signal if_stmt_956_branch_ack_1 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal addr_of_599_final_reg_req_0 : boolean;
  signal addr_of_599_final_reg_ack_0 : boolean;
  signal addr_of_599_final_reg_req_1 : boolean;
  signal addr_of_599_final_reg_ack_1 : boolean;
  signal type_cast_162_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_602_inst_req_0 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_602_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_602_inst_req_1 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_602_inst_ack_1 : boolean;
  signal if_stmt_956_branch_req_0 : boolean;
  signal type_cast_606_inst_req_0 : boolean;
  signal type_cast_606_inst_ack_0 : boolean;
  signal type_cast_606_inst_req_1 : boolean;
  signal type_cast_606_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_615_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_615_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_615_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_615_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 : boolean;
  signal ptr_deref_942_store_0_ack_1 : boolean;
  signal ptr_deref_942_store_0_req_1 : boolean;
  signal type_cast_619_inst_req_0 : boolean;
  signal type_cast_619_inst_ack_0 : boolean;
  signal type_cast_619_inst_req_1 : boolean;
  signal type_cast_619_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_633_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_633_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_633_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_633_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 : boolean;
  signal phi_stmt_189_req_1 : boolean;
  signal ptr_deref_942_store_0_ack_0 : boolean;
  signal ptr_deref_942_store_0_req_0 : boolean;
  signal type_cast_637_inst_req_0 : boolean;
  signal type_cast_637_inst_ack_0 : boolean;
  signal type_cast_637_inst_req_1 : boolean;
  signal type_cast_637_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_912_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_651_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_651_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_651_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_651_inst_ack_1 : boolean;
  signal type_cast_655_inst_req_0 : boolean;
  signal type_cast_655_inst_ack_0 : boolean;
  signal type_cast_655_inst_req_1 : boolean;
  signal type_cast_655_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_req_1 : boolean;
  signal phi_stmt_80_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_669_inst_ack_1 : boolean;
  signal type_cast_898_inst_ack_1 : boolean;
  signal type_cast_673_inst_req_0 : boolean;
  signal phi_stmt_73_ack_0 : boolean;
  signal type_cast_673_inst_ack_0 : boolean;
  signal type_cast_673_inst_req_1 : boolean;
  signal type_cast_673_inst_ack_1 : boolean;
  signal type_cast_898_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_687_inst_ack_1 : boolean;
  signal type_cast_691_inst_req_0 : boolean;
  signal type_cast_691_inst_ack_0 : boolean;
  signal type_cast_691_inst_req_1 : boolean;
  signal type_cast_691_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal ptr_deref_735_store_0_req_0 : boolean;
  signal ptr_deref_735_store_0_ack_0 : boolean;
  signal ptr_deref_735_store_0_req_1 : boolean;
  signal ptr_deref_735_store_0_ack_1 : boolean;
  signal if_stmt_749_branch_req_0 : boolean;
  signal if_stmt_749_branch_ack_1 : boolean;
  signal if_stmt_749_branch_ack_0 : boolean;
  signal type_cast_776_inst_req_0 : boolean;
  signal type_cast_776_inst_ack_0 : boolean;
  signal type_cast_776_inst_req_1 : boolean;
  signal type_cast_776_inst_ack_1 : boolean;
  signal array_obj_ref_805_index_offset_req_0 : boolean;
  signal array_obj_ref_805_index_offset_ack_0 : boolean;
  signal array_obj_ref_805_index_offset_req_1 : boolean;
  signal array_obj_ref_805_index_offset_ack_1 : boolean;
  signal addr_of_806_final_reg_req_0 : boolean;
  signal addr_of_806_final_reg_ack_0 : boolean;
  signal addr_of_806_final_reg_req_1 : boolean;
  signal addr_of_806_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_809_inst_ack_1 : boolean;
  signal type_cast_813_inst_req_0 : boolean;
  signal type_cast_813_inst_ack_0 : boolean;
  signal type_cast_813_inst_req_1 : boolean;
  signal type_cast_813_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_822_inst_ack_1 : boolean;
  signal type_cast_826_inst_req_0 : boolean;
  signal type_cast_826_inst_ack_0 : boolean;
  signal type_cast_826_inst_req_1 : boolean;
  signal type_cast_826_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_840_inst_ack_1 : boolean;
  signal type_cast_844_inst_req_0 : boolean;
  signal type_cast_844_inst_ack_0 : boolean;
  signal type_cast_844_inst_req_1 : boolean;
  signal type_cast_844_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 : boolean;
  signal type_cast_862_inst_req_0 : boolean;
  signal type_cast_862_inst_ack_0 : boolean;
  signal phi_stmt_270_req_0 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal phi_stmt_277_req_0 : boolean;
  signal type_cast_276_inst_req_0 : boolean;
  signal type_cast_276_inst_ack_0 : boolean;
  signal type_cast_276_inst_req_1 : boolean;
  signal type_cast_276_inst_ack_1 : boolean;
  signal phi_stmt_270_req_1 : boolean;
  signal type_cast_282_inst_req_0 : boolean;
  signal type_cast_282_inst_ack_0 : boolean;
  signal type_cast_282_inst_req_1 : boolean;
  signal type_cast_282_inst_ack_1 : boolean;
  signal phi_stmt_277_req_1 : boolean;
  signal phi_stmt_270_ack_0 : boolean;
  signal phi_stmt_277_ack_0 : boolean;
  signal type_cast_322_inst_req_0 : boolean;
  signal type_cast_322_inst_ack_0 : boolean;
  signal type_cast_322_inst_req_1 : boolean;
  signal type_cast_322_inst_ack_1 : boolean;
  signal phi_stmt_319_req_0 : boolean;
  signal phi_stmt_319_ack_0 : boolean;
  signal phi_stmt_586_req_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal phi_stmt_586_req_1 : boolean;
  signal phi_stmt_586_ack_0 : boolean;
  signal phi_stmt_793_req_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal phi_stmt_793_req_1 : boolean;
  signal phi_stmt_793_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(294 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(225);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/cr
      -- 
    rr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_47_store_0_req_1); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_62_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/rr
      -- 
    ca_106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_0); -- 
    rr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_38_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/ra
      -- 
    ra_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/ca
      -- 
    ca_120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/rr
      -- 
    rr_158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_47_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/ra
      -- 
    ra_159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/ca
      -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_start_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/cr
      -- 
    ra_179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/rr
      -- 
    ca_184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_62_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/ra
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/ca
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__exit__
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64__entry__
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_32/R_cmp208_65_place
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_else_link/$entry
      -- 
    branch_req_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_64_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	246 
    -- CP-element group 13: 	247 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/cr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$entry
      -- 
    if_choice_transition_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_160_inst_req_1); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_160_inst_req_0); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	233 
    -- CP-element group 14: 	234 
    -- CP-element group 14: 	235 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70__exit__
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    cr_2498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_1); -- 
    rr_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	241 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/ra
      -- 
    ra_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	241 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/ca
      -- 
    ca_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	241 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	33 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	241 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/req
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_102_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/ack
      -- 
    ack_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	241 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/rr
      -- 
    ack_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_105_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/ra
      -- 
    ra_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	241 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/ca
      -- 
    ca_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	241 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/rr
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_sample_start_
      -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_122_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(32) & testConfigure_CP_0_elements(241);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/ra
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_sample_completed_
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	241 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (12) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/merge_ack
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/rr
      -- 
    ca_375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    rr_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(25), ack => type_cast_126_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/ra
      -- 
    ra_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	241 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/ca
      -- 
    ca_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	241 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_update_start_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/cr
      -- 
    ra_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_137_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    cr_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(28), ack => RPIPE_ConvTranspose_input_pipe_137_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/rr
      -- 
    ca_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_137_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    rr_416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(29), ack => type_cast_141_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/ra
      -- 
    ra_417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_141_inst_ack_0, ack => testConfigure_CP_0_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	241 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/ca
      -- 
    ca_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_141_inst_ack_1, ack => testConfigure_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  delay-element  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	21 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_ptr_deref_122_delay
      -- 
    -- Element group testConfigure_CP_0_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  branch  join  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	17 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	27 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (10) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142__exit__
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143__entry__
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_dead_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/branch_req
      -- CP-element group 33: 	 branch_block_stmt_32/R_cmp_144_place
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_if_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_else_link/$entry
      -- 
    branch_req_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => if_stmt_143_branch_req_0); -- 
    testConfigure_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(27) & testConfigure_CP_0_elements(31);
      gj_testConfigure_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	226 
    -- CP-element group 34: 	227 
    -- CP-element group 34: 	229 
    -- CP-element group 34: 	230 
    -- CP-element group 34:  members (20) 
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/if_stmt_143_if_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/if_stmt_143_if_link/if_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/cr
      -- 
    if_choice_transition_436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_143_branch_ack_1, ack => testConfigure_CP_0_elements(34)); -- 
    rr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_76_inst_req_0); -- 
    cr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_76_inst_req_1); -- 
    rr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_83_inst_req_0); -- 
    cr_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_83_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	242 
    -- CP-element group 35: 	243 
    -- CP-element group 35:  members (12) 
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_143_else_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_143_else_link/else_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/cr
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    else_choice_transition_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_143_branch_ack_0, ack => testConfigure_CP_0_elements(35)); -- 
    cr_2534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => type_cast_153_inst_req_1); -- 
    rr_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => type_cast_153_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	253 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_171_store_0_ack_0, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  branch  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	253 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (15) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179__exit__
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180__entry__
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_dead_link/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/branch_req
      -- CP-element group 37: 	 branch_block_stmt_32/R_cmp14203_181_place
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_if_link/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_else_link/$entry
      -- 
    ca_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_171_store_0_ack_1, ack => testConfigure_CP_0_elements(37)); -- 
    branch_req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(37), ack => if_stmt_180_branch_req_0); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	260 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_32/if_stmt_180_if_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/if_stmt_180_if_link/if_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph200
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph200_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph200_PhiReq/$exit
      -- 
    if_choice_transition_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_180_branch_ack_1, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  merge  transition  place  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	257 
    -- CP-element group 39:  members (14) 
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186__exit__
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/dummy
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiReqMerge
      -- CP-element group 39: 	 branch_block_stmt_32/if_stmt_180_else_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/if_stmt_180_else_link/else_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$entry
      -- 
    else_choice_transition_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_180_branch_ack_0, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	259 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	259 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	59 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	259 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	59 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_sample_complete
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/ack
      -- 
    ack_557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_211_index_offset_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	259 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (11) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_offset_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/req
      -- 
    ack_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_211_index_offset_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    req_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(43), ack => addr_of_212_final_reg_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/ack
      -- 
    ack_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_212_final_reg_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	259 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (19) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/root_register_ack
      -- 
    ack_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_212_final_reg_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	259 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_update_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/cr
      -- 
    ra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_215_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    cr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(46), ack => RPIPE_ConvTranspose_input_pipe_215_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/rr
      -- 
    ca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_215_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    rr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(47), ack => type_cast_219_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/ra
      -- 
    ra_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => testConfigure_CP_0_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	259 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/ca
      -- 
    ca_605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/rr
      -- 
    rr_643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(50), ack => ptr_deref_222_store_0_req_0); -- 
    testConfigure_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(45) & testConfigure_CP_0_elements(49);
      gj_testConfigure_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	58 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/ra
      -- 
    ra_644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_store_0_ack_0, ack => testConfigure_CP_0_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	259 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	59 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/ca
      -- 
    ca_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_store_0_ack_1, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	259 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/rr
      -- 
    rr_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(53), ack => ptr_deref_239_load_0_req_0); -- 
    testConfigure_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(58) & testConfigure_CP_0_elements(259);
      gj_testConfigure_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/ra
      -- 
    ra_689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_0, ack => testConfigure_CP_0_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	259 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (12) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/merge_ack
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/rr
      -- 
    ca_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_1, ack => testConfigure_CP_0_elements(55)); -- 
    rr_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_243_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/ra
      -- 
    ra_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_0, ack => testConfigure_CP_0_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	259 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/ca
      -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_1, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  delay-element  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	53 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_ptr_deref_239_delay
      -- 
    -- Element group testConfigure_CP_0_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(51), ack => testConfigure_CP_0_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	41 
    -- CP-element group 59: 	42 
    -- CP-element group 59: 	52 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251__exit__
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252__entry__
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_32/R_cmp14_253_place
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_else_link/$entry
      -- 
    branch_req_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => if_stmt_252_branch_req_0); -- 
    testConfigure_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(41) & testConfigure_CP_0_elements(42) & testConfigure_CP_0_elements(52) & testConfigure_CP_0_elements(57);
      gj_testConfigure_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	254 
    -- CP-element group 60: 	255 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/cr
      -- CP-element group 60: 	 branch_block_stmt_32/if_stmt_252_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/if_stmt_252_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/$entry
      -- 
    if_choice_transition_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_1, ack => testConfigure_CP_0_elements(60)); -- 
    cr_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => type_cast_192_inst_req_1); -- 
    rr_2629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => type_cast_192_inst_req_0); -- 
    -- CP-element group 61:  merge  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	260 
    -- CP-element group 61:  members (13) 
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258__exit__
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph200x_xloopexit_bbx_xnph200
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/if_stmt_252_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/if_stmt_252_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph200x_xloopexit
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph200x_xloopexit_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph200x_xloopexit_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph200x_xloopexit_bbx_xnph200_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph200x_xloopexit_bbx_xnph200_PhiReq/$exit
      -- 
    else_choice_transition_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_0, ack => testConfigure_CP_0_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	260 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_update_start_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/cr
      -- 
    ra_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    cr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(62), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_1); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/rr
      -- 
    ca_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => type_cast_266_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/ra
      -- 
    ra_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	260 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	261 
    -- CP-element group 65: 	262 
    -- CP-element group 65: 	263 
    -- CP-element group 65:  members (17) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267__exit__
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/cr
      -- 
    ca_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    rr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(65), ack => type_cast_280_inst_req_0); -- 
    cr_2707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(65), ack => type_cast_280_inst_req_1); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	276 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/ack
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_sample_completed_
      -- 
    ack_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_287_final_reg_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	276 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (28) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_root_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_address_resized
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/base_resize_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/base_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/root_register_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/root_register_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/split_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/split_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/rr
      -- 
    ack_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_287_final_reg_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => ptr_deref_290_store_0_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/ra
      -- 
    ra_851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_290_store_0_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	276 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/ca
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_290_store_0_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	276 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_update_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/cr
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_0, ack => testConfigure_CP_0_elements(70)); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/rr
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_298_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/ra
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	276 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/ca
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_1, ack => testConfigure_CP_0_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311__exit__
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312__entry__
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_32/R_exitcond6_313_place
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_else_link/$entry
      -- 
    branch_req_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(74), ack => if_stmt_312_branch_req_0); -- 
    testConfigure_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(69) & testConfigure_CP_0_elements(73);
      gj_testConfigure_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	277 
    -- CP-element group 75: 	278 
    -- CP-element group 75:  members (12) 
      -- CP-element group 75: 	 branch_block_stmt_32/if_stmt_312_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/if_stmt_312_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/cr
      -- 
    if_choice_transition_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_312_branch_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(75), ack => type_cast_322_inst_req_0); -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(75), ack => type_cast_322_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	266 
    -- CP-element group 76: 	267 
    -- CP-element group 76: 	269 
    -- CP-element group 76: 	270 
    -- CP-element group 76:  members (20) 
      -- CP-element group 76: 	 branch_block_stmt_32/if_stmt_312_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/if_stmt_312_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/cr
      -- 
    else_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_312_branch_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_276_inst_req_0); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_276_inst_req_1); -- 
    rr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_282_inst_req_0); -- 
    cr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_282_inst_req_1); -- 
    -- CP-element group 77:  join  fork  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	280 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	80 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	86 
    -- CP-element group 77: 	90 
    -- CP-element group 77: 	91 
    -- CP-element group 77: 	93 
    -- CP-element group 77: 	97 
    -- CP-element group 77: 	98 
    -- CP-element group 77: 	100 
    -- CP-element group 77: 	101 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	104 
    -- CP-element group 77: 	105 
    -- CP-element group 77: 	106 
    -- CP-element group 77: 	108 
    -- CP-element group 77: 	109 
    -- CP-element group 77: 	110 
    -- CP-element group 77: 	112 
    -- CP-element group 77: 	113 
    -- CP-element group 77: 	114 
    -- CP-element group 77: 	116 
    -- CP-element group 77: 	117 
    -- CP-element group 77: 	118 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	122 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	125 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	128 
    -- CP-element group 77:  members (295) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/STORE_padding_324_Split/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/STORE_padding_324_Split/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/STORE_padding_324_Split/split_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/STORE_padding_324_Split/split_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Update/cr
      -- 
    cr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => STORE_padding_324_store_0_req_1); -- 
    rr_933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => STORE_padding_324_store_0_req_0); -- 
    rr_953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_0); -- 
    cr_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_332_inst_req_1); -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_343_store_0_req_1); -- 
    cr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_351_inst_req_1); -- 
    cr_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_362_store_0_req_1); -- 
    cr_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_370_inst_req_1); -- 
    cr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_381_store_0_req_1); -- 
    cr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_394_load_0_req_1); -- 
    rr_1212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_394_load_0_req_0); -- 
    cr_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_398_inst_req_1); -- 
    cr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_410_load_0_req_1); -- 
    rr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_410_load_0_req_0); -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_414_inst_req_1); -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_426_load_0_req_1); -- 
    rr_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_426_load_0_req_0); -- 
    cr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_430_inst_req_1); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_452_load_0_req_1); -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_452_load_0_req_0); -- 
    cr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_456_inst_req_1); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_468_load_0_req_1); -- 
    rr_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_468_load_0_req_0); -- 
    cr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_472_inst_req_1); -- 
    cr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_484_load_0_req_1); -- 
    rr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_484_load_0_req_0); -- 
    cr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_488_inst_req_1); -- 
    cr_1607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_500_load_0_req_1); -- 
    rr_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_500_load_0_req_0); -- 
    cr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_504_inst_req_1); -- 
    testConfigure_CP_0_elements(77) <= testConfigure_CP_0_elements(280);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Sample/word_access_start/word_0/ra
      -- 
    ra_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_324_store_0_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/STORE_padding_324_Update/word_access_complete/word_0/ca
      -- 
    ca_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_324_store_0_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_update_start_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Update/cr
      -- 
    ra_954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_0, ack => testConfigure_CP_0_elements(80)); -- 
    cr_958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	87 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_328_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Sample/rr
      -- 
    ca_959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_1, ack => testConfigure_CP_0_elements(81)); -- 
    rr_967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => type_cast_332_inst_req_0); -- 
    rr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Sample/ra
      -- 
    ra_968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_0, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_332_Update/ca
      -- 
    ca_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_1, ack => testConfigure_CP_0_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/ptr_deref_343_Split/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/ptr_deref_343_Split/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/ptr_deref_343_Split/split_req
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/ptr_deref_343_Split/split_ack
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/word_0/rr
      -- 
    rr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => ptr_deref_343_store_0_req_0); -- 
    testConfigure_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(83);
      gj_testConfigure_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	129 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Sample/word_access_start/word_0/ra
      -- 
    ra_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_store_0_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	77 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	131 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_Update/word_access_complete/word_0/ca
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_store_0_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_update_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Update/cr
      -- 
    ra_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_0, ack => testConfigure_CP_0_elements(87)); -- 
    cr_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	94 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_347_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- 
    ca_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_1, ack => testConfigure_CP_0_elements(88)); -- 
    rr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => type_cast_351_inst_req_0); -- 
    rr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Sample/ra
      -- 
    ra_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_0, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	77 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_351_Update/ca
      -- 
    ca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_1, ack => testConfigure_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	77 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	129 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/ptr_deref_362_Split/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/ptr_deref_362_Split/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/ptr_deref_362_Split/split_req
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/ptr_deref_362_Split/split_ack
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/word_0/rr
      -- 
    rr_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => ptr_deref_362_store_0_req_0); -- 
    testConfigure_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(90) & testConfigure_CP_0_elements(129);
      gj_testConfigure_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	130 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Sample/word_access_start/word_0/ra
      -- 
    ra_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_362_store_0_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	77 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	131 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_Update/word_access_complete/word_0/ca
      -- 
    ca_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_362_store_0_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	88 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => testConfigure_CP_0_elements(94)); -- 
    cr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_sample_start_
      -- 
    ca_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => testConfigure_CP_0_elements(95)); -- 
    rr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(95), ack => type_cast_370_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Sample/$exit
      -- 
    ra_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	77 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_370_update_completed_
      -- 
    ca_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	77 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	130 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/word_0/rr
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/ptr_deref_381_Split/split_ack
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/ptr_deref_381_Split/split_req
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/ptr_deref_381_Split/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/ptr_deref_381_Split/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/$entry
      -- 
    rr_1167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(98), ack => ptr_deref_381_store_0_req_0); -- 
    testConfigure_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(97) & testConfigure_CP_0_elements(130);
      gj_testConfigure_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Sample/$exit
      -- 
    ra_1168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_store_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	77 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	131 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_381_Update/$exit
      -- 
    ca_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_store_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	77 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_sample_completed_
      -- 
    ra_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (12) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/ptr_deref_394_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/ptr_deref_394_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/ptr_deref_394_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/ptr_deref_394_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_394_update_completed_
      -- 
    ca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    rr_1237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(102), ack => type_cast_398_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_sample_completed_
      -- 
    ra_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_398_inst_ack_0, ack => testConfigure_CP_0_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	77 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	131 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_398_update_completed_
      -- 
    ca_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_398_inst_ack_1, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	77 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/word_0/ra
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/word_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/word_access_start/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_sample_completed_
      -- 
    ra_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_410_load_0_ack_0, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	77 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (12) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/ptr_deref_410_Merge/merge_ack
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/ptr_deref_410_Merge/merge_req
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/ptr_deref_410_Merge/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/ptr_deref_410_Merge/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/word_0/ca
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/word_access_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_410_update_completed_
      -- 
    ca_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_410_load_0_ack_1, ack => testConfigure_CP_0_elements(106)); -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(106), ack => type_cast_414_inst_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_sample_completed_
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_414_inst_ack_0, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	77 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	131 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_414_update_completed_
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_414_inst_ack_1, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	77 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_sample_completed_
      -- 
    ra_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_0, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	77 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (12) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/ptr_deref_426_Merge/merge_ack
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/ptr_deref_426_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/ptr_deref_426_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/ptr_deref_426_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_426_update_completed_
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_1, ack => testConfigure_CP_0_elements(110)); -- 
    rr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(110), ack => type_cast_430_inst_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_sample_completed_
      -- 
    ra_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_0, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	77 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	131 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_430_update_completed_
      -- 
    ca_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_1, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	77 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/word_0/ra
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Sample/word_access_start/$exit
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_452_load_0_ack_0, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	77 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (12) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/ptr_deref_452_Merge/merge_ack
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/ptr_deref_452_Merge/merge_req
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/ptr_deref_452_Merge/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/ptr_deref_452_Merge/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/word_0/ca
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/word_access_complete/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_452_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Sample/$entry
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_452_load_0_ack_1, ack => testConfigure_CP_0_elements(114)); -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_456_inst_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Sample/$exit
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	77 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	131 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_456_Update/$exit
      -- 
    ca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	77 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/word_0/ra
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_sample_completed_
      -- 
    ra_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_0, ack => testConfigure_CP_0_elements(117)); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	77 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (12) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/ptr_deref_468_Merge/merge_ack
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/ptr_deref_468_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/ptr_deref_468_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_468_Update/ptr_deref_468_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Sample/$entry
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_1, ack => testConfigure_CP_0_elements(118)); -- 
    rr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_472_inst_req_0); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Sample/$exit
      -- 
    ra_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_0, ack => testConfigure_CP_0_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	131 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_472_update_completed_
      -- 
    ca_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/word_0/ra
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Sample/word_access_start/word_0/$exit
      -- 
    ra_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_484_load_0_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    -- CP-element group 122:  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	77 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (12) 
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/ptr_deref_484_Merge/merge_req
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/ptr_deref_484_Merge/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/ptr_deref_484_Merge/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/word_0/ca
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/word_0/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/word_access_complete/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_484_Update/ptr_deref_484_Merge/merge_ack
      -- 
    ca_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_484_load_0_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    rr_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(122), ack => type_cast_488_inst_req_0); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Sample/ra
      -- 
    ra_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_488_Update/ca
      -- 
    ca_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_1, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	77 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Sample/word_access_start/word_0/ra
      -- 
    ra_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_load_0_ack_0, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (12) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/word_access_complete/word_0/ca
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/ptr_deref_500_Merge/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/ptr_deref_500_Merge/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/ptr_deref_500_Merge/merge_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_500_Update/ptr_deref_500_Merge/merge_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Sample/rr
      -- 
    ca_1608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_load_0_ack_1, ack => testConfigure_CP_0_elements(126)); -- 
    rr_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(126), ack => type_cast_504_inst_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Sample/ra
      -- 
    ra_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => testConfigure_CP_0_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	77 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/type_cast_504_Update/ca
      -- 
    ca_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_1, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  transition  delay-element  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	85 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	91 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_343_ptr_deref_362_delay
      -- 
    -- Element group testConfigure_CP_0_elements(129) is a control-delay.
    cp_element_129_delay: control_delay_element  generic map(name => " 129_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(85), ack => testConfigure_CP_0_elements(129), clk => clk, reset =>reset);
    -- CP-element group 130:  transition  delay-element  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	92 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	98 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/ptr_deref_362_ptr_deref_381_delay
      -- 
    -- Element group testConfigure_CP_0_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(92), ack => testConfigure_CP_0_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  branch  join  transition  place  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: 	86 
    -- CP-element group 131: 	93 
    -- CP-element group 131: 	100 
    -- CP-element group 131: 	104 
    -- CP-element group 131: 	108 
    -- CP-element group 131: 	112 
    -- CP-element group 131: 	116 
    -- CP-element group 131: 	120 
    -- CP-element group 131: 	124 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (10) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526__exit__
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527__entry__
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_dead_link/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_eval_test/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_eval_test/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_eval_test/branch_req
      -- CP-element group 131: 	 branch_block_stmt_32/R_cmp71192_528_place
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_if_link/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_527_else_link/$entry
      -- 
    branch_req_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => if_stmt_527_branch_req_0); -- 
    testConfigure_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(79) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(104) & testConfigure_CP_0_elements(108) & testConfigure_CP_0_elements(112) & testConfigure_CP_0_elements(116) & testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(124) & testConfigure_CP_0_elements(128);
      gj_testConfigure_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	136 
    -- CP-element group 132: 	137 
    -- CP-element group 132:  members (18) 
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_548__exit__
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583__entry__
      -- CP-element group 132: 	 branch_block_stmt_32/if_stmt_527_if_link/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/if_stmt_527_if_link/if_choice_transition
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph194
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_update_start_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph194_PhiReq/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph194_PhiReq/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_548_PhiReqMerge
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_548_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_548_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_548_PhiAck/dummy
      -- 
    if_choice_transition_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_527_branch_ack_1, ack => testConfigure_CP_0_elements(132)); -- 
    rr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => type_cast_569_inst_req_0); -- 
    cr_1686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => type_cast_569_inst_req_1); -- 
    -- CP-element group 133:  transition  place  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	281 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_32/if_stmt_527_else_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/if_stmt_527_else_link/else_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond125x_xpreheader
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond125x_xpreheader_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond125x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_527_branch_ack_0, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	281 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	180 
    -- CP-element group 134: 	181 
    -- CP-element group 134:  members (18) 
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_755__exit__
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790__entry__
      -- CP-element group 134: 	 branch_block_stmt_32/if_stmt_542_if_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/if_stmt_542_if_link/if_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_bbx_xnph
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_update_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Update/cr
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_bbx_xnph_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_bbx_xnph_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_755_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_755_PhiAck/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_755_PhiAck/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_755_PhiAck/dummy
      -- 
    if_choice_transition_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_542_branch_ack_1, ack => testConfigure_CP_0_elements(134)); -- 
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => type_cast_776_inst_req_0); -- 
    cr_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => type_cast_776_inst_req_1); -- 
    -- CP-element group 135:  transition  place  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	281 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	294 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_542_else_link/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_542_else_link/else_choice_transition
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_forx_xend185
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_forx_xend185_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond125x_xpreheader_forx_xend185_PhiReq/$exit
      -- 
    else_choice_transition_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_542_branch_ack_0, ack => testConfigure_CP_0_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	132 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Sample/ra
      -- 
    ra_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  place  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	132 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	282 
    -- CP-element group 137:  members (9) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583__exit__
      -- CP-element group 137: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_554_to_assign_stmt_583/type_cast_569_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/$entry
      -- 
    ca_1687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	287 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	177 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_sample_complete
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Sample/ack
      -- 
    ack_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_598_index_offset_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    -- CP-element group 139:  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	287 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (11) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_offset_calculated
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_base_plus_offset/sum_rename_req
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_base_plus_offset/sum_rename_ack
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_request/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_request/req
      -- 
    ack_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_598_index_offset_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    req_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => addr_of_599_final_reg_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_request/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_request/ack
      -- 
    ack_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_599_final_reg_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	287 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	174 
    -- CP-element group 141:  members (19) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_complete/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_complete/ack
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_word_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_address_resized
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_addr_resize/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_addr_resize/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_addr_resize/base_resize_req
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_addr_resize/base_resize_ack
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_word_addrgen/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_word_addrgen/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_word_addrgen/root_register_req
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_word_addrgen/root_register_ack
      -- 
    ack_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_599_final_reg_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	287 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_update_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Update/cr
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_602_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_602_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Sample/rr
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_602_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    rr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => type_cast_606_inst_req_0); -- 
    rr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_615_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Sample/ra
      -- 
    ra_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	287 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	174 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Update/ca
      -- 
    ca_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_606_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_update_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Update/cr
      -- 
    ra_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_615_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    cr_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_615_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_615_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Sample/rr
      -- 
    ca_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_615_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    rr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => type_cast_619_inst_req_0); -- 
    rr_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_633_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Sample/ra
      -- 
    ra_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_619_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	287 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	174 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Update/ca
      -- 
    ca_1792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_619_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_update_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Update/cr
      -- 
    ra_1801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_633_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    cr_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_633_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_633_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Sample/rr
      -- 
    ca_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_633_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    rr_1814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => type_cast_637_inst_req_0); -- 
    rr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_651_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Sample/ra
      -- 
    ra_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_637_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	287 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	174 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Update/ca
      -- 
    ca_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_637_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_update_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Update/cr
      -- 
    ra_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_651_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_651_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_651_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Sample/rr
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_651_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    rr_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => type_cast_655_inst_req_0); -- 
    rr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_669_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Sample/ra
      -- 
    ra_1843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	287 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	174 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Update/ca
      -- 
    ca_1848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_655_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_update_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Update/cr
      -- 
    ra_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_669_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    cr_1861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(158), ack => RPIPE_ConvTranspose_input_pipe_669_inst_req_1); -- 
    -- CP-element group 159:  fork  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_669_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Sample/rr
      -- 
    ca_1862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_669_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    rr_1870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => type_cast_673_inst_req_0); -- 
    rr_1884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => RPIPE_ConvTranspose_input_pipe_687_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Sample/ra
      -- 
    ra_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	287 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	174 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Update/ca
      -- 
    ca_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_673_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	159 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (6) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_update_start_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Update/cr
      -- 
    ra_1885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_687_inst_ack_0, ack => testConfigure_CP_0_elements(162)); -- 
    cr_1889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(162), ack => RPIPE_ConvTranspose_input_pipe_687_inst_req_1); -- 
    -- CP-element group 163:  fork  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_687_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Sample/rr
      -- 
    ca_1890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_687_inst_ack_1, ack => testConfigure_CP_0_elements(163)); -- 
    rr_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(163), ack => type_cast_691_inst_req_0); -- 
    rr_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(163), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_0); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Sample/ra
      -- 
    ra_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_0, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	287 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	174 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Update/ca
      -- 
    ca_1904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_1, ack => testConfigure_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	163 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_update_start_
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Update/cr
      -- 
    ra_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_0, ack => testConfigure_CP_0_elements(166)); -- 
    cr_1917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(166), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_1); -- 
    -- CP-element group 167:  fork  transition  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: 	170 
    -- CP-element group 167:  members (9) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_705_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Sample/rr
      -- 
    ca_1918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_1, ack => testConfigure_CP_0_elements(167)); -- 
    rr_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_709_inst_req_0); -- 
    rr_1940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_0); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Sample/ra
      -- 
    ra_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	287 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	174 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Update/ca
      -- 
    ca_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	167 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_update_start_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Update/cr
      -- 
    ra_1941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    cr_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(170), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_1); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_723_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Sample/rr
      -- 
    ca_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    rr_1954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(171), ack => type_cast_727_inst_req_0); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Sample/ra
      -- 
    ra_1955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	287 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Update/ca
      -- 
    ca_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	141 
    -- CP-element group 174: 	145 
    -- CP-element group 174: 	149 
    -- CP-element group 174: 	153 
    -- CP-element group 174: 	157 
    -- CP-element group 174: 	161 
    -- CP-element group 174: 	165 
    -- CP-element group 174: 	169 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/ptr_deref_735_Split/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/ptr_deref_735_Split/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/ptr_deref_735_Split/split_req
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/ptr_deref_735_Split/split_ack
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/word_0/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/word_0/rr
      -- 
    rr_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => ptr_deref_735_store_0_req_0); -- 
    testConfigure_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(145) & testConfigure_CP_0_elements(149) & testConfigure_CP_0_elements(153) & testConfigure_CP_0_elements(157) & testConfigure_CP_0_elements(161) & testConfigure_CP_0_elements(165) & testConfigure_CP_0_elements(169) & testConfigure_CP_0_elements(173);
      gj_testConfigure_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (5) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/word_0/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Sample/word_access_start/word_0/ra
      -- 
    ra_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_735_store_0_ack_0, ack => testConfigure_CP_0_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	287 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (5) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/word_0/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/word_0/ca
      -- 
    ca_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_735_store_0_ack_1, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  branch  join  transition  place  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	138 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (10) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748__exit__
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749__entry__
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_dead_link/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_eval_test/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_eval_test/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_eval_test/branch_req
      -- CP-element group 177: 	 branch_block_stmt_32/R_exitcond_750_place
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_if_link/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_749_else_link/$entry
      -- 
    branch_req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(177), ack => if_stmt_749_branch_req_0); -- 
    testConfigure_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(138) & testConfigure_CP_0_elements(176);
      gj_testConfigure_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  merge  transition  place  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	281 
    -- CP-element group 178:  members (13) 
      -- CP-element group 178: 	 branch_block_stmt_32/merge_stmt_533__exit__
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xcond125x_xpreheaderx_xloopexit_forx_xcond125x_xpreheader
      -- CP-element group 178: 	 branch_block_stmt_32/if_stmt_749_if_link/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/if_stmt_749_if_link/if_choice_transition
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xbody73_forx_xcond125x_xpreheaderx_xloopexit
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xbody73_forx_xcond125x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xbody73_forx_xcond125x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/merge_stmt_533_PhiReqMerge
      -- CP-element group 178: 	 branch_block_stmt_32/merge_stmt_533_PhiAck/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/merge_stmt_533_PhiAck/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/merge_stmt_533_PhiAck/dummy
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xcond125x_xpreheaderx_xloopexit_forx_xcond125x_xpreheader_PhiReq/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/forx_xcond125x_xpreheaderx_xloopexit_forx_xcond125x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_2023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_749_branch_ack_1, ack => testConfigure_CP_0_elements(178)); -- 
    -- CP-element group 179:  fork  transition  place  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	283 
    -- CP-element group 179: 	284 
    -- CP-element group 179:  members (12) 
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_749_else_link/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_749_else_link/else_choice_transition
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_749_branch_ack_0, ack => testConfigure_CP_0_elements(179)); -- 
    rr_2864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_592_inst_req_0); -- 
    cr_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_592_inst_req_1); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	134 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Sample/ra
      -- 
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  place  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	134 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	288 
    -- CP-element group 181:  members (9) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790__exit__
      -- CP-element group 181: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_761_to_assign_stmt_790/type_cast_776_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/$entry
      -- 
    ca_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	293 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	221 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_sample_complete
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Sample/ack
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_805_index_offset_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	293 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (11) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_root_address_calculated
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_offset_calculated
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Update/ack
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_base_plus_offset/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_base_plus_offset/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_base_plus_offset/sum_rename_req
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_base_plus_offset/sum_rename_ack
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_request/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_request/req
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_805_index_offset_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    req_2089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => addr_of_806_final_reg_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_request/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_request/ack
      -- 
    ack_2090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_806_final_reg_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  fork  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	293 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	218 
    -- CP-element group 185:  members (19) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_word_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_root_address_calculated
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_address_resized
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_addr_resize/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_word_addrgen/root_register_ack
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_word_addrgen/root_register_req
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_word_addrgen/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_word_addrgen/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_plus_offset/sum_rename_ack
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_plus_offset/sum_rename_req
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_plus_offset/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_plus_offset/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_addr_resize/base_resize_ack
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_addr_resize/base_resize_req
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_base_addr_resize/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_complete/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_complete/ack
      -- 
    ack_2095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_806_final_reg_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	293 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_update_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Update/cr
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_809_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_809_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Sample/rr
      -- 
    ca_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_809_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_813_inst_req_0); -- 
    rr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_822_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Sample/ra
      -- 
    ra_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	293 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	218 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Update/ca
      -- 
    ca_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_update_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Update/cr
      -- 
    ra_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_822_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_822_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_822_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Sample/rr
      -- 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_822_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_826_inst_req_0); -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_840_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Sample/ra
      -- 
    ra_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	293 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	218 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Update/ca
      -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_update_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Update/cr
      -- 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_840_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_840_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_840_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Sample/rr
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_840_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_844_inst_req_0); -- 
    rr_2187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Sample/ra
      -- 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	293 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	218 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Update/ca
      -- 
    ca_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_844_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_update_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Update/cr
      -- 
    ra_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_858_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_858_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Sample/rr
      -- 
    ca_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_858_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_862_inst_req_0); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Sample/ra
      -- 
    ra_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	293 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	218 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_update_completed_
      -- 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_862_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_update_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Update/cr
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Update/$entry
      -- 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_876_inst_req_1); -- 
    -- CP-element group 203:  fork  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203: 	206 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_876_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_sample_start_
      -- 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_876_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_880_inst_req_0); -- 
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Sample/ra
      -- 
    ra_2230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	293 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	218 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Update/ca
      -- 
    ca_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	203 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Update/cr
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Sample/ra
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_update_start_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_sample_completed_
      -- 
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_0, ack => testConfigure_CP_0_elements(206)); -- 
    cr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => RPIPE_ConvTranspose_input_pipe_894_inst_req_1); -- 
    -- CP-element group 207:  fork  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	210 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Update/ca
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_894_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_sample_start_
      -- 
    ca_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_894_inst_ack_1, ack => testConfigure_CP_0_elements(207)); -- 
    rr_2257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => type_cast_898_inst_req_0); -- 
    rr_2271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_0); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Sample/ra
      -- 
    ra_2258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_0, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	293 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	218 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Update/ca
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Update/$exit
      -- 
    ca_2263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_1, ack => testConfigure_CP_0_elements(209)); -- 
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	207 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (6) 
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Sample/ra
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Sample/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_update_start_
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_sample_completed_
      -- 
    ra_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_0, ack => testConfigure_CP_0_elements(210)); -- 
    cr_2276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(210), ack => RPIPE_ConvTranspose_input_pipe_912_inst_req_1); -- 
    -- CP-element group 211:  fork  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211: 	214 
    -- CP-element group 211:  members (9) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Update/ca
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_Update/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_912_update_completed_
      -- 
    ca_2277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_912_inst_ack_1, ack => testConfigure_CP_0_elements(211)); -- 
    rr_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_916_inst_req_0); -- 
    rr_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => RPIPE_ConvTranspose_input_pipe_930_inst_req_0); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_sample_completed_
      -- 
    ra_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	293 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_update_completed_
      -- 
    ca_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	211 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_update_start_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Sample/ra
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Update/cr
      -- 
    ra_2300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_930_inst_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    cr_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(214), ack => RPIPE_ConvTranspose_input_pipe_930_inst_req_1); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Update/ca
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_930_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Sample/rr
      -- 
    ca_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_930_inst_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    rr_2313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(215), ack => type_cast_934_inst_req_0); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Sample/ra
      -- 
    ra_2314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_0, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	293 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Update/ca
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Update/$exit
      -- 
    ca_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_934_inst_ack_1, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	185 
    -- CP-element group 218: 	189 
    -- CP-element group 218: 	193 
    -- CP-element group 218: 	197 
    -- CP-element group 218: 	201 
    -- CP-element group 218: 	205 
    -- CP-element group 218: 	209 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (9) 
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/word_0/rr
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/word_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/ptr_deref_942_Split/split_ack
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/ptr_deref_942_Split/split_req
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/ptr_deref_942_Split/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/ptr_deref_942_Split/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/$entry
      -- 
    rr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(218), ack => ptr_deref_942_store_0_req_0); -- 
    testConfigure_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205) & testConfigure_CP_0_elements(209) & testConfigure_CP_0_elements(213) & testConfigure_CP_0_elements(217);
      gj_testConfigure_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/word_0/ra
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/word_0/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/word_access_start/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Sample/$exit
      -- 
    ra_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_store_0_ack_0, ack => testConfigure_CP_0_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	293 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/word_0/ca
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/word_0/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/$exit
      -- 
    ca_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_store_0_ack_1, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  branch  join  transition  place  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	182 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (10) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956__entry__
      -- CP-element group 221: 	 branch_block_stmt_32/R_exitcond5_957_place
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_else_link/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_if_link/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_eval_test/branch_req
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_eval_test/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_eval_test/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/if_stmt_956_dead_link/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/$exit
      -- 
    branch_req_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(221), ack => if_stmt_956_branch_req_0); -- 
    testConfigure_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(182) & testConfigure_CP_0_elements(220);
      gj_testConfigure_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  merge  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	294 
    -- CP-element group 222:  members (13) 
      -- CP-element group 222: 	 branch_block_stmt_32/merge_stmt_962__exit__
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xend185x_xloopexit_forx_xend185
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbody131_forx_xend185x_xloopexit
      -- CP-element group 222: 	 branch_block_stmt_32/if_stmt_956_if_link/if_choice_transition
      -- CP-element group 222: 	 branch_block_stmt_32/if_stmt_956_if_link/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbody131_forx_xend185x_xloopexit_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbody131_forx_xend185x_xloopexit_PhiReq/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/merge_stmt_962_PhiReqMerge
      -- CP-element group 222: 	 branch_block_stmt_32/merge_stmt_962_PhiAck/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/merge_stmt_962_PhiAck/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/merge_stmt_962_PhiAck/dummy
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xend185x_xloopexit_forx_xend185_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xend185x_xloopexit_forx_xend185_PhiReq/$exit
      -- 
    if_choice_transition_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_1, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  fork  transition  place  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	289 
    -- CP-element group 223: 	290 
    -- CP-element group 223:  members (12) 
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131
      -- CP-element group 223: 	 branch_block_stmt_32/if_stmt_956_else_link/else_choice_transition
      -- CP-element group 223: 	 branch_block_stmt_32/if_stmt_956_else_link/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/rr
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_0, ack => testConfigure_CP_0_elements(223)); -- 
    rr_2918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(223), ack => type_cast_799_inst_req_0); -- 
    cr_2923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(223), ack => type_cast_799_inst_req_1); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	294 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Sample/ra
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_sample_completed_
      -- 
    ra_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => testConfigure_CP_0_elements(224)); -- 
    -- CP-element group 225:  transition  place  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	294 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (16) 
      -- CP-element group 225: 	 $exit
      -- CP-element group 225: 	 branch_block_stmt_32/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_968__exit__
      -- CP-element group 225: 	 branch_block_stmt_32/return__
      -- CP-element group 225: 	 branch_block_stmt_32/merge_stmt_970__exit__
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Update/ca
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_968/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/merge_stmt_970_PhiReqMerge
      -- CP-element group 225: 	 branch_block_stmt_32/merge_stmt_970_PhiAck/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/merge_stmt_970_PhiAck/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/merge_stmt_970_PhiAck/dummy
      -- 
    ca_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	34 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/ra
      -- 
    ra_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => testConfigure_CP_0_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	34 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (2) 
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/ca
      -- 
    ca_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => testConfigure_CP_0_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	232 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$exit
      -- 
    phi_stmt_73_req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(228), ack => phi_stmt_73_req_0); -- 
    testConfigure_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(226) & testConfigure_CP_0_elements(227);
      gj_testConfigure_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	34 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (2) 
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/ra
      -- 
    ra_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => testConfigure_CP_0_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	34 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (2) 
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/ca
      -- 
    ca_2465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  join  transition  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => phi_stmt_80_req_0); -- 
    testConfigure_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(229) & testConfigure_CP_0_elements(230);
      gj_testConfigure_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  join  transition  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	228 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	238 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(228) & testConfigure_CP_0_elements(231);
      gj_testConfigure_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  output  delay-element  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	14 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	237 
    -- CP-element group 233:  members (4) 
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_79_konst_delay_trans
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- 
    phi_stmt_73_req_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(233), ack => phi_stmt_73_req_1); -- 
    -- Element group testConfigure_CP_0_elements(233) is a control-delay.
    cp_element_233_delay: control_delay_element  generic map(name => " 233_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(233), clk => clk, reset =>reset);
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	14 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/ra
      -- 
    ra_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	14 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/ca
      -- 
    ca_2499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_80_req_1); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	233 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(233) & testConfigure_CP_0_elements(236);
      gj_testConfigure_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  merge  fork  transition  place  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	232 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_32/merge_stmt_72_PhiReqMerge
      -- CP-element group 238: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(238) <= OrReduce(testConfigure_CP_0_elements(232) & testConfigure_CP_0_elements(237));
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (1) 
      -- CP-element group 239: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_73_ack
      -- 
    phi_stmt_73_ack_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_73_ack_0, ack => testConfigure_CP_0_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_80_ack
      -- 
    phi_stmt_80_ack_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_80_ack_0, ack => testConfigure_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  fork  transition  place  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	15 
    -- CP-element group 241: 	16 
    -- CP-element group 241: 	17 
    -- CP-element group 241: 	18 
    -- CP-element group 241: 	20 
    -- CP-element group 241: 	22 
    -- CP-element group 241: 	23 
    -- CP-element group 241: 	25 
    -- CP-element group 241: 	27 
    -- CP-element group 241: 	28 
    -- CP-element group 241: 	31 
    -- CP-element group 241:  members (64) 
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_72__exit__
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142__entry__
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/root_register_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/root_register_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/rr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resized_1
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scaled_1
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_computed_1
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/index_resize_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/index_resize_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/scale_rename_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/scale_rename_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_update_start
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/cr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_root_address_calculated
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_address_resized
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/base_resize_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/base_resize_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/sum_rename_req
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/sum_rename_ack
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/cr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/rr
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/cr
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$exit
      -- 
    rr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_95_inst_req_0); -- 
    cr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_95_inst_req_1); -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => array_obj_ref_101_index_offset_req_0); -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => array_obj_ref_101_index_offset_req_1); -- 
    req_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => addr_of_102_final_reg_req_1); -- 
    cr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => ptr_deref_105_store_0_req_1); -- 
    cr_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => ptr_deref_122_load_0_req_1); -- 
    cr_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_126_inst_req_1); -- 
    rr_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => RPIPE_ConvTranspose_input_pipe_137_inst_req_0); -- 
    cr_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_141_inst_req_1); -- 
    testConfigure_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(239) & testConfigure_CP_0_elements(240);
      gj_testConfigure_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	35 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$exit
      -- 
    ra_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	35 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/ca
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$exit
      -- 
    ca_2535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  place  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (8) 
      -- CP-element group 244: 	 branch_block_stmt_32/merge_stmt_149_PhiReqMerge
      -- CP-element group 244: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$entry
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- 
    phi_stmt_150_req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_150_req_0); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	249 
    -- CP-element group 245: 	250 
    -- CP-element group 245:  members (13) 
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/cr
      -- CP-element group 245: 	 branch_block_stmt_32/merge_stmt_149__exit__
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/phi_stmt_150_ack
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/rr
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/$entry
      -- 
    phi_stmt_150_ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => testConfigure_CP_0_elements(245)); -- 
    cr_2591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(245), ack => type_cast_162_inst_req_1); -- 
    rr_2586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(245), ack => type_cast_162_inst_req_0); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	13 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/ra
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_0, ack => testConfigure_CP_0_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	13 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (2) 
      -- CP-element group 247: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/ca
      -- CP-element group 247: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/$exit
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_1, ack => testConfigure_CP_0_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	252 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_req
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_157_req_2567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_157_req_2567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(248), ack => phi_stmt_157_req_0); -- 
    testConfigure_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(246) & testConfigure_CP_0_elements(247);
      gj_testConfigure_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	245 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (2) 
      -- CP-element group 249: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/ra
      -- CP-element group 249: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/$exit
      -- 
    ra_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_0, ack => testConfigure_CP_0_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	245 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/ca
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/$exit
      -- 
    ca_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_1, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  join  transition  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_req
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/$exit
      -- 
    phi_stmt_157_req_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_157_req_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(251), ack => phi_stmt_157_req_1); -- 
    testConfigure_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(249) & testConfigure_CP_0_elements(250);
      gj_testConfigure_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  merge  transition  place  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	248 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (2) 
      -- CP-element group 252: 	 branch_block_stmt_32/merge_stmt_156_PhiReqMerge
      -- CP-element group 252: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(252) <= OrReduce(testConfigure_CP_0_elements(248) & testConfigure_CP_0_elements(251));
    -- CP-element group 253:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	36 
    -- CP-element group 253: 	37 
    -- CP-element group 253:  members (35) 
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_156__exit__
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179__entry__
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/phi_stmt_157_ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_address_calculated
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_address_calculated
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_root_address_calculated
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_address_resized
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/base_resize_req
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/base_resize_ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/sum_rename_req
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/sum_rename_ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/root_register_req
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/root_register_ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/split_req
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/split_ack
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/rr
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/cr
      -- 
    phi_stmt_157_ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_157_ack_0, ack => testConfigure_CP_0_elements(253)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => ptr_deref_171_store_0_req_0); -- 
    cr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => ptr_deref_171_store_0_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	60 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/ra
      -- CP-element group 254: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/$exit
      -- 
    ra_2630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_0, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	60 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/ca
      -- CP-element group 255: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/$exit
      -- 
    ca_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_1, ack => testConfigure_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_req
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/$exit
      -- 
    phi_stmt_189_req_2636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_189_req_2636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => phi_stmt_189_req_0); -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(254) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  output  delay-element  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	39 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_req
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_195_konst_delay_trans
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$exit
      -- 
    phi_stmt_189_req_2647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_189_req_2647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(257), ack => phi_stmt_189_req_1); -- 
    -- Element group testConfigure_CP_0_elements(257) is a control-delay.
    cp_element_257_delay: control_delay_element  generic map(name => " 257_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(39), ack => testConfigure_CP_0_elements(257), clk => clk, reset =>reset);
    -- CP-element group 258:  merge  transition  place  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/merge_stmt_188_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(258) <= OrReduce(testConfigure_CP_0_elements(256) & testConfigure_CP_0_elements(257));
    -- CP-element group 259:  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	40 
    -- CP-element group 259: 	41 
    -- CP-element group 259: 	42 
    -- CP-element group 259: 	43 
    -- CP-element group 259: 	45 
    -- CP-element group 259: 	46 
    -- CP-element group 259: 	49 
    -- CP-element group 259: 	52 
    -- CP-element group 259: 	53 
    -- CP-element group 259: 	55 
    -- CP-element group 259: 	57 
    -- CP-element group 259:  members (65) 
      -- CP-element group 259: 	 branch_block_stmt_32/merge_stmt_188__exit__
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251__entry__
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resized_1
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scaled_1
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_computed_1
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/index_resize_req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/index_resize_ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/scale_rename_req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/scale_rename_ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_update_start
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/cr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_address_calculated
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_address_calculated
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_root_address_calculated
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_address_resized
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/base_resize_req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/base_resize_ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/sum_rename_req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/sum_rename_ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/root_register_req
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/root_register_ack
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/cr
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/cr
      -- CP-element group 259: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/phi_stmt_189_ack
      -- CP-element group 259: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/$exit
      -- 
    phi_stmt_189_ack_2652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_189_ack_0, ack => testConfigure_CP_0_elements(259)); -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => type_cast_205_inst_req_0); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => type_cast_205_inst_req_1); -- 
    req_556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => array_obj_ref_211_index_offset_req_0); -- 
    req_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => array_obj_ref_211_index_offset_req_1); -- 
    req_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => addr_of_212_final_reg_req_1); -- 
    rr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => RPIPE_ConvTranspose_input_pipe_215_inst_req_0); -- 
    cr_604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => type_cast_219_inst_req_1); -- 
    cr_654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => ptr_deref_222_store_0_req_1); -- 
    cr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => ptr_deref_239_load_0_req_1); -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => type_cast_243_inst_req_1); -- 
    -- CP-element group 260:  merge  fork  transition  place  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	38 
    -- CP-element group 260: 	61 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	62 
    -- CP-element group 260: 	65 
    -- CP-element group 260:  members (13) 
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_260__exit__
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267__entry__
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_update_start_
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/cr
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_260_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/dummy
      -- 
    rr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_0); -- 
    cr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => type_cast_266_inst_req_1); -- 
    testConfigure_CP_0_elements(260) <= OrReduce(testConfigure_CP_0_elements(38) & testConfigure_CP_0_elements(61));
    -- CP-element group 261:  transition  output  delay-element  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	65 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	265 
    -- CP-element group 261:  members (4) 
      -- CP-element group 261: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_274_konst_delay_trans
      -- CP-element group 261: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_req
      -- 
    phi_stmt_270_req_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_270_req_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => phi_stmt_270_req_0); -- 
    -- Element group testConfigure_CP_0_elements(261) is a control-delay.
    cp_element_261_delay: control_delay_element  generic map(name => " 261_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(65), ack => testConfigure_CP_0_elements(261), clk => clk, reset =>reset);
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	65 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/ra
      -- 
    ra_2703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	65 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/ca
      -- 
    ca_2708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (5) 
      -- CP-element group 264: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_req
      -- 
    phi_stmt_277_req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_277_req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => phi_stmt_277_req_0); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	261 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	273 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_32/bbx_xnph200_forx_xbody30_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(261) & testConfigure_CP_0_elements(264);
      gj_testConfigure_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	76 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/ra
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_0, ack => testConfigure_CP_0_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	76 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (2) 
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/ca
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_1, ack => testConfigure_CP_0_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	272 
    -- CP-element group 268:  members (5) 
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_req
      -- 
    phi_stmt_270_req_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_270_req_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => phi_stmt_270_req_1); -- 
    testConfigure_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(266) & testConfigure_CP_0_elements(267);
      gj_testConfigure_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	76 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/ra
      -- 
    ra_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_0, ack => testConfigure_CP_0_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	76 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/ca
      -- 
    ca_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_1, ack => testConfigure_CP_0_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (5) 
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_req
      -- 
    phi_stmt_277_req_2758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_277_req_2758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => phi_stmt_277_req_1); -- 
    testConfigure_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(269) & testConfigure_CP_0_elements(270);
      gj_testConfigure_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  join  transition  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	268 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (1) 
      -- CP-element group 272: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(268) & testConfigure_CP_0_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  merge  fork  transition  place  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	265 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_32/merge_stmt_269_PhiReqMerge
      -- CP-element group 273: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(273) <= OrReduce(testConfigure_CP_0_elements(265) & testConfigure_CP_0_elements(272));
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/phi_stmt_270_ack
      -- 
    phi_stmt_270_ack_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_270_ack_0, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/phi_stmt_277_ack
      -- 
    phi_stmt_277_ack_2764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_277_ack_0, ack => testConfigure_CP_0_elements(275)); -- 
    -- CP-element group 276:  join  fork  transition  place  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	66 
    -- CP-element group 276: 	67 
    -- CP-element group 276: 	69 
    -- CP-element group 276: 	70 
    -- CP-element group 276: 	73 
    -- CP-element group 276:  members (42) 
      -- CP-element group 276: 	 branch_block_stmt_32/merge_stmt_269__exit__
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311__entry__
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/scale_rename_req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/scale_rename_ack
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/ack
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/sum_rename_req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/sum_rename_ack
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_update_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_root_address_calculated
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_offset_calculated
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resized_0
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scaled_0
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_computed_0
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/index_resize_req
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/index_resize_ack
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_update_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/cr
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/rr
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_update_start_
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/cr
      -- CP-element group 276: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/$exit
      -- 
    req_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => addr_of_287_final_reg_req_0); -- 
    req_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => addr_of_287_final_reg_req_1); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => ptr_deref_290_store_0_req_1); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_0); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => type_cast_298_inst_req_1); -- 
    testConfigure_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(274) & testConfigure_CP_0_elements(275);
      gj_testConfigure_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	75 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	75 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_1, ack => testConfigure_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  place  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (8) 
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_req
      -- CP-element group 279: 	 branch_block_stmt_32/merge_stmt_318_PhiReqMerge
      -- CP-element group 279: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/$entry
      -- 
    phi_stmt_319_req_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_319_req_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => phi_stmt_319_req_0); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  merge  transition  place  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	77 
    -- CP-element group 280:  members (4) 
      -- CP-element group 280: 	 branch_block_stmt_32/merge_stmt_318__exit__
      -- CP-element group 280: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_526__entry__
      -- CP-element group 280: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/phi_stmt_319_ack
      -- 
    phi_stmt_319_ack_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_319_ack_0, ack => testConfigure_CP_0_elements(280)); -- 
    -- CP-element group 281:  merge  branch  transition  place  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	133 
    -- CP-element group 281: 	178 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	134 
    -- CP-element group 281: 	135 
    -- CP-element group 281:  members (17) 
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_535__exit__
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_541__entry__
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_541__exit__
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542__entry__
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_541/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/assign_stmt_541/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_dead_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_eval_test/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_eval_test/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_eval_test/branch_req
      -- CP-element group 281: 	 branch_block_stmt_32/R_cmp129189_543_place
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_if_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/if_stmt_542_else_link/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_535_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_535_PhiAck/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_535_PhiAck/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_535_PhiAck/dummy
      -- 
    branch_req_1659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => if_stmt_542_branch_req_0); -- 
    testConfigure_CP_0_elements(281) <= OrReduce(testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(178));
    -- CP-element group 282:  transition  output  delay-element  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	137 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	286 
    -- CP-element group 282:  members (5) 
      -- CP-element group 282: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_590_konst_delay_trans
      -- CP-element group 282: 	 branch_block_stmt_32/bbx_xnph194_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_req
      -- 
    phi_stmt_586_req_2845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_586_req_2845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(282), ack => phi_stmt_586_req_0); -- 
    -- Element group testConfigure_CP_0_elements(282) is a control-delay.
    cp_element_282_delay: control_delay_element  generic map(name => " 282_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(137), ack => testConfigure_CP_0_elements(282), clk => clk, reset =>reset);
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	179 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Sample/ra
      -- 
    ra_2865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => testConfigure_CP_0_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	179 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/Update/ca
      -- 
    ca_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => testConfigure_CP_0_elements(284)); -- 
    -- CP-element group 285:  join  transition  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_sources/type_cast_592/SplitProtocol/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody73_forx_xbody73_PhiReq/phi_stmt_586/phi_stmt_586_req
      -- 
    phi_stmt_586_req_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_586_req_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(285), ack => phi_stmt_586_req_1); -- 
    testConfigure_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(283) & testConfigure_CP_0_elements(284);
      gj_testConfigure_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  merge  transition  place  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	282 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_32/merge_stmt_585_PhiReqMerge
      -- CP-element group 286: 	 branch_block_stmt_32/merge_stmt_585_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(286) <= OrReduce(testConfigure_CP_0_elements(282) & testConfigure_CP_0_elements(285));
    -- CP-element group 287:  fork  transition  place  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	138 
    -- CP-element group 287: 	139 
    -- CP-element group 287: 	141 
    -- CP-element group 287: 	142 
    -- CP-element group 287: 	145 
    -- CP-element group 287: 	149 
    -- CP-element group 287: 	153 
    -- CP-element group 287: 	157 
    -- CP-element group 287: 	161 
    -- CP-element group 287: 	165 
    -- CP-element group 287: 	169 
    -- CP-element group 287: 	173 
    -- CP-element group 287: 	176 
    -- CP-element group 287:  members (56) 
      -- CP-element group 287: 	 branch_block_stmt_32/merge_stmt_585__exit__
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748__entry__
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_resized_1
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_scaled_1
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_computed_1
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_resize_1/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_resize_1/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_resize_1/index_resize_req
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_resize_1/index_resize_ack
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_scale_1/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_scale_1/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_scale_1/scale_rename_req
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_index_scale_1/scale_rename_ack
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_update_start
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Sample/req
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/array_obj_ref_598_final_index_sum_regn_Update/req
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_complete/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/addr_of_599_complete/req
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/RPIPE_ConvTranspose_input_pipe_602_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_606_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_619_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_637_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_655_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_673_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_691_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_709_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/type_cast_727_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/word_0/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/assign_stmt_600_to_assign_stmt_748/ptr_deref_735_Update/word_access_complete/word_0/cr
      -- CP-element group 287: 	 branch_block_stmt_32/merge_stmt_585_PhiAck/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/merge_stmt_585_PhiAck/phi_stmt_586_ack
      -- 
    phi_stmt_586_ack_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_586_ack_0, ack => testConfigure_CP_0_elements(287)); -- 
    req_1715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => array_obj_ref_598_index_offset_req_0); -- 
    req_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => array_obj_ref_598_index_offset_req_1); -- 
    req_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => addr_of_599_final_reg_req_1); -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => RPIPE_ConvTranspose_input_pipe_602_inst_req_0); -- 
    cr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_606_inst_req_1); -- 
    cr_1791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_619_inst_req_1); -- 
    cr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_637_inst_req_1); -- 
    cr_1847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_655_inst_req_1); -- 
    cr_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_673_inst_req_1); -- 
    cr_1903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_691_inst_req_1); -- 
    cr_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_709_inst_req_1); -- 
    cr_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => type_cast_727_inst_req_1); -- 
    cr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => ptr_deref_735_store_0_req_1); -- 
    -- CP-element group 288:  transition  output  delay-element  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	181 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	292 
    -- CP-element group 288:  members (5) 
      -- CP-element group 288: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_797_konst_delay_trans
      -- CP-element group 288: 	 branch_block_stmt_32/bbx_xnph_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_req
      -- 
    phi_stmt_793_req_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_793_req_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(288), ack => phi_stmt_793_req_0); -- 
    -- Element group testConfigure_CP_0_elements(288) is a control-delay.
    cp_element_288_delay: control_delay_element  generic map(name => " 288_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(181), ack => testConfigure_CP_0_elements(288), clk => clk, reset =>reset);
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	223 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/ra
      -- 
    ra_2919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => testConfigure_CP_0_elements(289)); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	223 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (2) 
      -- CP-element group 290: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/ca
      -- 
    ca_2924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => testConfigure_CP_0_elements(290)); -- 
    -- CP-element group 291:  join  transition  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody131_forx_xbody131_PhiReq/phi_stmt_793/phi_stmt_793_req
      -- 
    phi_stmt_793_req_2925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_793_req_2925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(291), ack => phi_stmt_793_req_1); -- 
    testConfigure_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(289) & testConfigure_CP_0_elements(290);
      gj_testConfigure_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  merge  transition  place  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	288 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_32/merge_stmt_792_PhiReqMerge
      -- CP-element group 292: 	 branch_block_stmt_32/merge_stmt_792_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(292) <= OrReduce(testConfigure_CP_0_elements(288) & testConfigure_CP_0_elements(291));
    -- CP-element group 293:  fork  transition  place  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	182 
    -- CP-element group 293: 	183 
    -- CP-element group 293: 	185 
    -- CP-element group 293: 	186 
    -- CP-element group 293: 	189 
    -- CP-element group 293: 	193 
    -- CP-element group 293: 	197 
    -- CP-element group 293: 	201 
    -- CP-element group 293: 	205 
    -- CP-element group 293: 	209 
    -- CP-element group 293: 	213 
    -- CP-element group 293: 	217 
    -- CP-element group 293: 	220 
    -- CP-element group 293:  members (56) 
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/merge_stmt_792__exit__
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955__entry__
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_880_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_934_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_916_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/word_0/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/word_0/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/word_access_complete/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/ptr_deref_942_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_898_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_resized_1
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_scaled_1
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_computed_1
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_resize_1/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_resize_1/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_resize_1/index_resize_req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_resize_1/index_resize_ack
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_scale_1/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_scale_1/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_scale_1/scale_rename_req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_index_scale_1/scale_rename_ack
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_update_start
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/array_obj_ref_805_final_index_sum_regn_Update/req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_complete/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/addr_of_806_complete/req
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/RPIPE_ConvTranspose_input_pipe_809_Sample/rr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_813_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_826_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_844_Update/cr
      -- CP-element group 293: 	 branch_block_stmt_32/assign_stmt_807_to_assign_stmt_955/type_cast_862_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/merge_stmt_792_PhiAck/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/merge_stmt_792_PhiAck/phi_stmt_793_ack
      -- 
    phi_stmt_793_ack_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_793_ack_0, ack => testConfigure_CP_0_elements(293)); -- 
    cr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_934_inst_req_1); -- 
    cr_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_916_inst_req_1); -- 
    cr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_880_inst_req_1); -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_862_inst_req_1); -- 
    cr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => ptr_deref_942_store_0_req_1); -- 
    cr_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_898_inst_req_1); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => array_obj_ref_805_index_offset_req_0); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => array_obj_ref_805_index_offset_req_1); -- 
    req_2094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => addr_of_806_final_reg_req_1); -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => RPIPE_ConvTranspose_input_pipe_809_inst_req_0); -- 
    cr_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_813_inst_req_1); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_826_inst_req_1); -- 
    cr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => type_cast_844_inst_req_1); -- 
    -- CP-element group 294:  merge  fork  transition  place  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	135 
    -- CP-element group 294: 	222 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	224 
    -- CP-element group 294: 	225 
    -- CP-element group 294:  members (13) 
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_964__exit__
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968__entry__
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Update/cr
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Sample/rr
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_update_start_
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/type_cast_967_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_32/assign_stmt_968/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_964_PhiReqMerge
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_964_PhiAck/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_964_PhiAck/$exit
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_964_PhiAck/dummy
      -- 
    cr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(294), ack => type_cast_967_inst_req_1); -- 
    rr_2399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(294), ack => type_cast_967_inst_req_0); -- 
    testConfigure_CP_0_elements(294) <= OrReduce(testConfigure_CP_0_elements(135) & testConfigure_CP_0_elements(222));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar226_597_resized : std_logic_vector(13 downto 0);
    signal R_indvar226_597_scaled : std_logic_vector(13 downto 0);
    signal R_indvar241_285_resized : std_logic_vector(0 downto 0);
    signal R_indvar241_285_scaled : std_logic_vector(0 downto 0);
    signal R_indvar244_210_resized : std_logic_vector(6 downto 0);
    signal R_indvar244_210_scaled : std_logic_vector(6 downto 0);
    signal R_indvar249_100_resized : std_logic_vector(6 downto 0);
    signal R_indvar249_100_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_804_resized : std_logic_vector(10 downto 0);
    signal R_indvar_804_scaled : std_logic_vector(10 downto 0);
    signal STORE_padding_324_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_324_word_address_0 : std_logic_vector(0 downto 0);
    signal add104_697 : std_logic_vector(63 downto 0);
    signal add110_715 : std_logic_vector(63 downto 0);
    signal add116_733 : std_logic_vector(63 downto 0);
    signal add141_832 : std_logic_vector(63 downto 0);
    signal add147_850 : std_logic_vector(63 downto 0);
    signal add153_868 : std_logic_vector(63 downto 0);
    signal add159_886 : std_logic_vector(63 downto 0);
    signal add165_904 : std_logic_vector(63 downto 0);
    signal add171_922 : std_logic_vector(63 downto 0);
    signal add177_940 : std_logic_vector(63 downto 0);
    signal add86_643 : std_logic_vector(63 downto 0);
    signal add92_661 : std_logic_vector(63 downto 0);
    signal add98_679 : std_logic_vector(63 downto 0);
    signal add_625 : std_logic_vector(63 downto 0);
    signal array_obj_ref_101_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_286_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_598_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_598_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_598_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_598_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_598_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_598_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_805_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_805_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_805_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_805_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_805_root_address : std_logic_vector(10 downto 0);
    signal arrayidx120_600 : std_logic_vector(31 downto 0);
    signal arrayidx181_807 : std_logic_vector(31 downto 0);
    signal arrayidx21_213 : std_logic_vector(31 downto 0);
    signal arrayidx35_288 : std_logic_vector(31 downto 0);
    signal arrayidx_103 : std_logic_vector(31 downto 0);
    signal call101_688 : std_logic_vector(7 downto 0);
    signal call107_706 : std_logic_vector(7 downto 0);
    signal call113_724 : std_logic_vector(7 downto 0);
    signal call134_810 : std_logic_vector(7 downto 0);
    signal call138_823 : std_logic_vector(7 downto 0);
    signal call144_841 : std_logic_vector(7 downto 0);
    signal call150_859 : std_logic_vector(7 downto 0);
    signal call156_877 : std_logic_vector(7 downto 0);
    signal call162_895 : std_logic_vector(7 downto 0);
    signal call168_913 : std_logic_vector(7 downto 0);
    signal call174_931 : std_logic_vector(7 downto 0);
    signal call17_216 : std_logic_vector(7 downto 0);
    signal call31196_263 : std_logic_vector(7 downto 0);
    signal call31_295 : std_logic_vector(7 downto 0);
    signal call4209_59 : std_logic_vector(7 downto 0);
    signal call42_329 : std_logic_vector(7 downto 0);
    signal call44_348 : std_logic_vector(7 downto 0);
    signal call46_367 : std_logic_vector(7 downto 0);
    signal call4_138 : std_logic_vector(7 downto 0);
    signal call75_603 : std_logic_vector(7 downto 0);
    signal call78_616 : std_logic_vector(7 downto 0);
    signal call83_634 : std_logic_vector(7 downto 0);
    signal call89_652 : std_logic_vector(7 downto 0);
    signal call95_670 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp129189_541 : std_logic_vector(0 downto 0);
    signal cmp14203_179 : std_logic_vector(0 downto 0);
    signal cmp14_251 : std_logic_vector(0 downto 0);
    signal cmp208_56 : std_logic_vector(0 downto 0);
    signal cmp71192_526 : std_logic_vector(0 downto 0);
    signal cmp_135 : std_logic_vector(0 downto 0);
    signal conv103_692 : std_logic_vector(63 downto 0);
    signal conv109_710 : std_logic_vector(63 downto 0);
    signal conv115_728 : std_logic_vector(63 downto 0);
    signal conv135_814 : std_logic_vector(63 downto 0);
    signal conv13_244 : std_logic_vector(31 downto 0);
    signal conv140_827 : std_logic_vector(63 downto 0);
    signal conv146_845 : std_logic_vector(63 downto 0);
    signal conv152_863 : std_logic_vector(63 downto 0);
    signal conv158_881 : std_logic_vector(63 downto 0);
    signal conv164_899 : std_logic_vector(63 downto 0);
    signal conv170_917 : std_logic_vector(63 downto 0);
    signal conv176_935 : std_logic_vector(63 downto 0);
    signal conv18_220 : std_logic_vector(15 downto 0);
    signal conv2_127 : std_logic_vector(31 downto 0);
    signal conv32197_267 : std_logic_vector(15 downto 0);
    signal conv32199_277 : std_logic_vector(15 downto 0);
    signal conv32_299 : std_logic_vector(15 downto 0);
    signal conv32x_xlcssa_319 : std_logic_vector(15 downto 0);
    signal conv43_333 : std_logic_vector(15 downto 0);
    signal conv45_352 : std_logic_vector(15 downto 0);
    signal conv47_371 : std_logic_vector(15 downto 0);
    signal conv50_399 : std_logic_vector(31 downto 0);
    signal conv5210_63 : std_logic_vector(15 downto 0);
    signal conv5212_80 : std_logic_vector(15 downto 0);
    signal conv52_415 : std_logic_vector(31 downto 0);
    signal conv54_431 : std_logic_vector(31 downto 0);
    signal conv58_457 : std_logic_vector(31 downto 0);
    signal conv5_142 : std_logic_vector(15 downto 0);
    signal conv5x_xlcssa1_150 : std_logic_vector(15 downto 0);
    signal conv5x_xlcssa_157 : std_logic_vector(15 downto 0);
    signal conv60_473 : std_logic_vector(31 downto 0);
    signal conv63_489 : std_logic_vector(31 downto 0);
    signal conv66_505 : std_logic_vector(31 downto 0);
    signal conv76_607 : std_logic_vector(63 downto 0);
    signal conv80_620 : std_logic_vector(63 downto 0);
    signal conv85_638 : std_logic_vector(63 downto 0);
    signal conv91_656 : std_logic_vector(63 downto 0);
    signal conv97_674 : std_logic_vector(63 downto 0);
    signal conv_39 : std_logic_vector(15 downto 0);
    signal exitcond5_955 : std_logic_vector(0 downto 0);
    signal exitcond6_311 : std_logic_vector(0 downto 0);
    signal exitcond_748 : std_logic_vector(0 downto 0);
    signal iNsTr_13_119 : std_logic_vector(31 downto 0);
    signal iNsTr_1_45 : std_logic_vector(31 downto 0);
    signal iNsTr_21_236 : std_logic_vector(31 downto 0);
    signal iNsTr_26_341 : std_logic_vector(31 downto 0);
    signal iNsTr_29_360 : std_logic_vector(31 downto 0);
    signal iNsTr_32_379 : std_logic_vector(31 downto 0);
    signal iNsTr_34_391 : std_logic_vector(31 downto 0);
    signal iNsTr_35_407 : std_logic_vector(31 downto 0);
    signal iNsTr_36_423 : std_logic_vector(31 downto 0);
    signal iNsTr_37_449 : std_logic_vector(31 downto 0);
    signal iNsTr_38_465 : std_logic_vector(31 downto 0);
    signal iNsTr_39_481 : std_logic_vector(31 downto 0);
    signal iNsTr_40_497 : std_logic_vector(31 downto 0);
    signal iNsTr_43_570 : std_logic_vector(63 downto 0);
    signal iNsTr_56_777 : std_logic_vector(63 downto 0);
    signal iNsTr_5_169 : std_logic_vector(31 downto 0);
    signal inc24_206 : std_logic_vector(31 downto 0);
    signal inc_96 : std_logic_vector(31 downto 0);
    signal indvar226_586 : std_logic_vector(63 downto 0);
    signal indvar241_270 : std_logic_vector(63 downto 0);
    signal indvar244_189 : std_logic_vector(63 downto 0);
    signal indvar249_73 : std_logic_vector(63 downto 0);
    signal indvar_793 : std_logic_vector(63 downto 0);
    signal indvarx_xnext227_743 : std_logic_vector(63 downto 0);
    signal indvarx_xnext242_305 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_950 : std_logic_vector(63 downto 0);
    signal mul55_441 : std_logic_vector(31 downto 0);
    signal mul61_510 : std_logic_vector(31 downto 0);
    signal mul64_515 : std_logic_vector(31 downto 0);
    signal mul67_520 : std_logic_vector(31 downto 0);
    signal mul_436 : std_logic_vector(31 downto 0);
    signal ptr_deref_105_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_105_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_105_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_105_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_122_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_171_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_171_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_171_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_171_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_171_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_171_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_222_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_222_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_222_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_222_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_222_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_222_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_239_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_239_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_239_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_239_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_239_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_290_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_290_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_290_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_290_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_290_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_290_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_343_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_343_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_343_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_343_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_362_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_362_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_362_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_362_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_362_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_362_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_381_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_381_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_394_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_410_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_410_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_410_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_410_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_410_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_426_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_452_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_452_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_452_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_452_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_452_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_468_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_47_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_47_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_484_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_484_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_484_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_484_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_484_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_500_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_500_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_500_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_500_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_500_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_735_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_735_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_735_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_735_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_735_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_735_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_942_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_942_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_942_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_942_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_942_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_942_word_offset_0 : std_logic_vector(10 downto 0);
    signal shl100_685 : std_logic_vector(63 downto 0);
    signal shl106_703 : std_logic_vector(63 downto 0);
    signal shl112_721 : std_logic_vector(63 downto 0);
    signal shl137_820 : std_logic_vector(63 downto 0);
    signal shl143_838 : std_logic_vector(63 downto 0);
    signal shl149_856 : std_logic_vector(63 downto 0);
    signal shl155_874 : std_logic_vector(63 downto 0);
    signal shl161_892 : std_logic_vector(63 downto 0);
    signal shl167_910 : std_logic_vector(63 downto 0);
    signal shl173_928 : std_logic_vector(63 downto 0);
    signal shl82_631 : std_logic_vector(63 downto 0);
    signal shl88_649 : std_logic_vector(63 downto 0);
    signal shl94_667 : std_logic_vector(63 downto 0);
    signal shl_613 : std_logic_vector(63 downto 0);
    signal tmp12_240 : std_logic_vector(15 downto 0);
    signal tmp1_123 : std_logic_vector(15 downto 0);
    signal tmp221_761 : std_logic_vector(31 downto 0);
    signal tmp221x_xop_773 : std_logic_vector(31 downto 0);
    signal tmp222_767 : std_logic_vector(0 downto 0);
    signal tmp225_790 : std_logic_vector(63 downto 0);
    signal tmp233_554 : std_logic_vector(31 downto 0);
    signal tmp233x_xop_566 : std_logic_vector(31 downto 0);
    signal tmp234_560 : std_logic_vector(0 downto 0);
    signal tmp238_583 : std_logic_vector(63 downto 0);
    signal tmp246_230 : std_logic_vector(63 downto 0);
    signal tmp251_113 : std_logic_vector(63 downto 0);
    signal tmp3_202 : std_logic_vector(63 downto 0);
    signal tmp49_395 : std_logic_vector(15 downto 0);
    signal tmp51_411 : std_logic_vector(15 downto 0);
    signal tmp53_427 : std_logic_vector(15 downto 0);
    signal tmp57_453 : std_logic_vector(15 downto 0);
    signal tmp59_469 : std_logic_vector(15 downto 0);
    signal tmp62_485 : std_logic_vector(15 downto 0);
    signal tmp65_501 : std_logic_vector(15 downto 0);
    signal tmp_92 : std_logic_vector(63 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_131_wire : std_logic_vector(31 downto 0);
    signal type_cast_133_wire : std_logic_vector(31 downto 0);
    signal type_cast_153_wire : std_logic_vector(15 downto 0);
    signal type_cast_160_wire : std_logic_vector(15 downto 0);
    signal type_cast_162_wire : std_logic_vector(15 downto 0);
    signal type_cast_177_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_192_wire : std_logic_vector(63 downto 0);
    signal type_cast_195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_200_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_228_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_247_wire : std_logic_vector(31 downto 0);
    signal type_cast_249_wire : std_logic_vector(31 downto 0);
    signal type_cast_274_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_276_wire : std_logic_vector(63 downto 0);
    signal type_cast_280_wire : std_logic_vector(15 downto 0);
    signal type_cast_282_wire : std_logic_vector(15 downto 0);
    signal type_cast_303_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_309_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_322_wire : std_logic_vector(15 downto 0);
    signal type_cast_524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_539_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_53_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_552_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_564_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_574_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_581_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_592_wire : std_logic_vector(63 downto 0);
    signal type_cast_611_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_629_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_683_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_741_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_76_wire : std_logic_vector(63 downto 0);
    signal type_cast_771_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_799_wire : std_logic_vector(63 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_83_wire : std_logic_vector(15 downto 0);
    signal type_cast_854_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire : std_logic_vector(15 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop253_576 : std_logic_vector(63 downto 0);
    signal xx_xop_783 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_324_word_address_0 <= "0";
    array_obj_ref_101_constant_part_of_offset <= "0000011";
    array_obj_ref_101_offset_scale_factor_0 <= "1000000";
    array_obj_ref_101_offset_scale_factor_1 <= "0000001";
    array_obj_ref_101_resized_base_address <= "0000000";
    array_obj_ref_211_constant_part_of_offset <= "0000011";
    array_obj_ref_211_offset_scale_factor_0 <= "1000000";
    array_obj_ref_211_offset_scale_factor_1 <= "0000001";
    array_obj_ref_211_resized_base_address <= "0000000";
    array_obj_ref_286_offset_scale_factor_0 <= "1";
    array_obj_ref_286_resized_base_address <= "0";
    array_obj_ref_598_constant_part_of_offset <= "00000000000000";
    array_obj_ref_598_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_598_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_598_resized_base_address <= "00000000000000";
    array_obj_ref_805_constant_part_of_offset <= "00000010001";
    array_obj_ref_805_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_805_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_805_resized_base_address <= "00000000000";
    iNsTr_13_119 <= "00000000000000000000000000000010";
    iNsTr_1_45 <= "00000000000000000000000000000010";
    iNsTr_21_236 <= "00000000000000000000000000000010";
    iNsTr_26_341 <= "00000000000000000000000000000011";
    iNsTr_29_360 <= "00000000000000000000000000000100";
    iNsTr_32_379 <= "00000000000000000000000000000101";
    iNsTr_34_391 <= "00000000000000000000000000000011";
    iNsTr_35_407 <= "00000000000000000000000000000100";
    iNsTr_36_423 <= "00000000000000000000000000000101";
    iNsTr_37_449 <= "00000000000000000000000000000011";
    iNsTr_38_465 <= "00000000000000000000000000000100";
    iNsTr_39_481 <= "00000000000000000000000000000101";
    iNsTr_40_497 <= "00000000000000000000000000000110";
    iNsTr_5_169 <= "00000000000000000000000000000010";
    ptr_deref_105_word_offset_0 <= "0000000";
    ptr_deref_122_word_offset_0 <= "0000000";
    ptr_deref_171_word_offset_0 <= "0000000";
    ptr_deref_222_word_offset_0 <= "0000000";
    ptr_deref_239_word_offset_0 <= "0000000";
    ptr_deref_290_word_offset_0 <= "0";
    ptr_deref_343_word_offset_0 <= "0000000";
    ptr_deref_362_word_offset_0 <= "0000000";
    ptr_deref_381_word_offset_0 <= "0000000";
    ptr_deref_394_word_offset_0 <= "0000000";
    ptr_deref_410_word_offset_0 <= "0000000";
    ptr_deref_426_word_offset_0 <= "0000000";
    ptr_deref_452_word_offset_0 <= "0000000";
    ptr_deref_468_word_offset_0 <= "0000000";
    ptr_deref_47_word_offset_0 <= "0000000";
    ptr_deref_484_word_offset_0 <= "0000000";
    ptr_deref_500_word_offset_0 <= "0000000";
    ptr_deref_735_word_offset_0 <= "00000000000000";
    ptr_deref_942_word_offset_0 <= "00000000000";
    type_cast_111_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_177_wire_constant <= "0000000000000000";
    type_cast_195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_200_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_228_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_274_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_309_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_524_wire_constant <= "00000000000000000000000000000011";
    type_cast_539_wire_constant <= "00000000000000000000000000000011";
    type_cast_53_wire_constant <= "00000000";
    type_cast_552_wire_constant <= "00000000000000000000000000000010";
    type_cast_558_wire_constant <= "00000000000000000000000000000001";
    type_cast_564_wire_constant <= "11111111111111111111111111111111";
    type_cast_574_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_581_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_590_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_611_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_629_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_647_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_665_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_683_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_741_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_759_wire_constant <= "00000000000000000000000000000010";
    type_cast_765_wire_constant <= "00000000000000000000000000000001";
    type_cast_771_wire_constant <= "11111111111111111111111111111111";
    type_cast_781_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_79_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_836_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_854_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_90_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire;
      req(0) <= phi_stmt_150_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => conv5x_xlcssa1_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    phi_stmt_157: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_160_wire & type_cast_162_wire;
      req <= phi_stmt_157_req_0 & phi_stmt_157_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_157",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_157_ack_0,
          idata => idata,
          odata => conv5x_xlcssa_157,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_157
    phi_stmt_189: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_192_wire & type_cast_195_wire_constant;
      req <= phi_stmt_189_req_0 & phi_stmt_189_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_189",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_189_ack_0,
          idata => idata,
          odata => indvar244_189,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_189
    phi_stmt_270: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_274_wire_constant & type_cast_276_wire;
      req <= phi_stmt_270_req_0 & phi_stmt_270_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_270",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_270_ack_0,
          idata => idata,
          odata => indvar241_270,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_270
    phi_stmt_277: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_280_wire & type_cast_282_wire;
      req <= phi_stmt_277_req_0 & phi_stmt_277_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_277",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_277_ack_0,
          idata => idata,
          odata => conv32199_277,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_277
    phi_stmt_319: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_322_wire;
      req(0) <= phi_stmt_319_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_319",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_319_ack_0,
          idata => idata,
          odata => conv32x_xlcssa_319,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_319
    phi_stmt_586: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_590_wire_constant & type_cast_592_wire;
      req <= phi_stmt_586_req_0 & phi_stmt_586_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_586",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_586_ack_0,
          idata => idata,
          odata => indvar226_586,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_586
    phi_stmt_73: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire & type_cast_79_wire_constant;
      req <= phi_stmt_73_req_0 & phi_stmt_73_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_73",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_73_ack_0,
          idata => idata,
          odata => indvar249_73,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_73
    phi_stmt_793: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_797_wire_constant & type_cast_799_wire;
      req <= phi_stmt_793_req_0 & phi_stmt_793_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_793",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_793_ack_0,
          idata => idata,
          odata => indvar_793,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_793
    phi_stmt_80: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_83_wire & type_cast_85_wire;
      req <= phi_stmt_80_req_0 & phi_stmt_80_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_80",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_80_ack_0,
          idata => idata,
          odata => conv5212_80,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_80
    -- flow-through select operator MUX_582_inst
    tmp238_583 <= xx_xop253_576 when (tmp234_560(0) /=  '0') else type_cast_581_wire_constant;
    -- flow-through select operator MUX_789_inst
    tmp225_790 <= xx_xop_783 when (tmp222_767(0) /=  '0') else type_cast_788_wire_constant;
    addr_of_102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_102_final_reg_req_0;
      addr_of_102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_102_final_reg_req_1;
      addr_of_102_final_reg_ack_1<= rack(0);
      addr_of_102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_212_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_212_final_reg_req_0;
      addr_of_212_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_212_final_reg_req_1;
      addr_of_212_final_reg_ack_1<= rack(0);
      addr_of_212_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_212_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_211_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx21_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_287_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_287_final_reg_req_0;
      addr_of_287_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_287_final_reg_req_1;
      addr_of_287_final_reg_ack_1<= rack(0);
      addr_of_287_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_287_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_286_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx35_288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_599_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_599_final_reg_req_0;
      addr_of_599_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_599_final_reg_req_1;
      addr_of_599_final_reg_ack_1<= rack(0);
      addr_of_599_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_599_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_598_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx120_600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_806_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_806_final_reg_req_0;
      addr_of_806_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_806_final_reg_req_1;
      addr_of_806_final_reg_ack_1<= rack(0);
      addr_of_806_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_806_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_805_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx181_807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_131_inst
    process(inc_96) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc_96(31 downto 0);
      type_cast_131_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_133_inst
    process(conv2_127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv2_127(31 downto 0);
      type_cast_133_wire <= tmp_var; -- 
    end process;
    type_cast_141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_141_inst_req_0;
      type_cast_141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_141_inst_req_1;
      type_cast_141_inst_ack_1<= rack(0);
      type_cast_141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5_142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_160_inst_req_0;
      type_cast_160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_160_inst_req_1;
      type_cast_160_inst_ack_1<= rack(0);
      type_cast_160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5210_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_160_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_162_inst_req_0;
      type_cast_162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_162_inst_req_1;
      type_cast_162_inst_ack_1<= rack(0);
      type_cast_162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5x_xlcssa1_150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_162_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_192_inst_req_0;
      type_cast_192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_192_inst_req_1;
      type_cast_192_inst_ack_1<= rack(0);
      type_cast_192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp246_230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_192_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc24_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call17_216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_243_inst_req_0;
      type_cast_243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_243_inst_req_1;
      type_cast_243_inst_ack_1<= rack(0);
      type_cast_243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_247_inst
    process(inc24_206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc24_206(31 downto 0);
      type_cast_247_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_249_inst
    process(conv13_244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv13_244(31 downto 0);
      type_cast_249_wire <= tmp_var; -- 
    end process;
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31196_263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32197_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_276_inst_req_0;
      type_cast_276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_276_inst_req_1;
      type_cast_276_inst_ack_1<= rack(0);
      type_cast_276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext242_305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_276_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32197_267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_280_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_282_inst_req_0;
      type_cast_282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_282_inst_req_1;
      type_cast_282_inst_ack_1<= rack(0);
      type_cast_282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_282_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_298_inst_req_0;
      type_cast_298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_298_inst_req_1;
      type_cast_298_inst_ack_1<= rack(0);
      type_cast_298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_295,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_322_inst_req_0;
      type_cast_322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_322_inst_req_1;
      type_cast_322_inst_ack_1<= rack(0);
      type_cast_322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_322_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_332_inst_req_0;
      type_cast_332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_332_inst_req_1;
      type_cast_332_inst_ack_1<= rack(0);
      type_cast_332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_351_inst_req_0;
      type_cast_351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_351_inst_req_1;
      type_cast_351_inst_ack_1<= rack(0);
      type_cast_351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_398_inst_req_0;
      type_cast_398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_398_inst_req_1;
      type_cast_398_inst_ack_1<= rack(0);
      type_cast_398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp49_395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_414_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_414_inst_req_0;
      type_cast_414_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_414_inst_req_1;
      type_cast_414_inst_ack_1<= rack(0);
      type_cast_414_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_414_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp51_411,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_430_inst_req_0;
      type_cast_430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_430_inst_req_1;
      type_cast_430_inst_ack_1<= rack(0);
      type_cast_430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp53_427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp57_453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_472_inst_req_0;
      type_cast_472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_472_inst_req_1;
      type_cast_472_inst_ack_1<= rack(0);
      type_cast_472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp59_469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_488_inst_req_0;
      type_cast_488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_488_inst_req_1;
      type_cast_488_inst_ack_1<= rack(0);
      type_cast_488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp62_485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_504_inst_req_1;
      type_cast_504_inst_ack_1<= rack(0);
      type_cast_504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp65_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_569_inst_req_0;
      type_cast_569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_569_inst_req_1;
      type_cast_569_inst_ack_1<= rack(0);
      type_cast_569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp233x_xop_566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_43_570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext227_743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_592_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_606_inst_req_0;
      type_cast_606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_606_inst_req_1;
      type_cast_606_inst_ack_1<= rack(0);
      type_cast_606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call75_603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_619_inst_req_0;
      type_cast_619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_619_inst_req_1;
      type_cast_619_inst_ack_1<= rack(0);
      type_cast_619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call78_616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_62_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_62_inst_req_0;
      type_cast_62_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_62_inst_req_1;
      type_cast_62_inst_ack_1<= rack(0);
      type_cast_62_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_62_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4209_59,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5210_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_637_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_637_inst_req_0;
      type_cast_637_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_637_inst_req_1;
      type_cast_637_inst_ack_1<= rack(0);
      type_cast_637_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_637_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call83_634,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_638,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_655_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_655_inst_req_0;
      type_cast_655_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_655_inst_req_1;
      type_cast_655_inst_ack_1<= rack(0);
      type_cast_655_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_655_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_652,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_673_inst_req_0;
      type_cast_673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_673_inst_req_1;
      type_cast_673_inst_ack_1<= rack(0);
      type_cast_673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_691_inst_req_0;
      type_cast_691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_691_inst_req_1;
      type_cast_691_inst_ack_1<= rack(0);
      type_cast_691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_688,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call113_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp251_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_76_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_776_inst_req_0;
      type_cast_776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_776_inst_req_1;
      type_cast_776_inst_ack_1<= rack(0);
      type_cast_776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp221x_xop_773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_56_777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_813_inst_req_0;
      type_cast_813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_813_inst_req_1;
      type_cast_813_inst_ack_1<= rack(0);
      type_cast_813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_826_inst_req_0;
      type_cast_826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_826_inst_req_1;
      type_cast_826_inst_ack_1<= rack(0);
      type_cast_826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv140_827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_83_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_844_inst_req_0;
      type_cast_844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_844_inst_req_1;
      type_cast_844_inst_ack_1<= rack(0);
      type_cast_844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call144_841,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5210_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_85_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_862_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_862_inst_req_0;
      type_cast_862_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_862_inst_req_1;
      type_cast_862_inst_ack_1<= rack(0);
      type_cast_862_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_862_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call150_859,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv152_863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_880_inst_req_0;
      type_cast_880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_880_inst_req_1;
      type_cast_880_inst_ack_1<= rack(0);
      type_cast_880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call156_877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_898_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_898_inst_req_0;
      type_cast_898_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_898_inst_req_1;
      type_cast_898_inst_ack_1<= rack(0);
      type_cast_898_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_898_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call162_895,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv164_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_934_inst_req_0;
      type_cast_934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_934_inst_req_1;
      type_cast_934_inst_ack_1<= rack(0);
      type_cast_934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_935,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul55_441,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_324_gather_scatter
    process(conv32x_xlcssa_319) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv32x_xlcssa_319;
      ov(15 downto 0) := iv;
      STORE_padding_324_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_rename
    process(R_indvar249_100_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar249_100_resized;
      ov(6 downto 0) := iv;
      R_indvar249_100_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_resize
    process(indvar249_73) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar249_73;
      ov := iv(6 downto 0);
      R_indvar249_100_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_root_address_inst
    process(array_obj_ref_101_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_101_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_index_1_rename
    process(R_indvar244_210_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar244_210_resized;
      ov(6 downto 0) := iv;
      R_indvar244_210_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_index_1_resize
    process(indvar244_189) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar244_189;
      ov := iv(6 downto 0);
      R_indvar244_210_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_root_address_inst
    process(array_obj_ref_211_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_211_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_211_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_0_rename
    process(R_indvar241_285_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar241_285_resized;
      ov(0 downto 0) := iv;
      R_indvar241_285_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_0_resize
    process(indvar241_270) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar241_270;
      ov := iv(0 downto 0);
      R_indvar241_285_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_offset
    process(R_indvar241_285_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar241_285_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_286_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_root_address_inst
    process(array_obj_ref_286_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_286_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_286_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_598_index_1_rename
    process(R_indvar226_597_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar226_597_resized;
      ov(13 downto 0) := iv;
      R_indvar226_597_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_598_index_1_resize
    process(indvar226_586) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar226_586;
      ov := iv(13 downto 0);
      R_indvar226_597_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_598_root_address_inst
    process(array_obj_ref_598_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_598_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_598_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_index_1_rename
    process(R_indvar_804_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_804_resized;
      ov(10 downto 0) := iv;
      R_indvar_804_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_index_1_resize
    process(indvar_793) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_793;
      ov := iv(10 downto 0);
      R_indvar_804_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_root_address_inst
    process(array_obj_ref_805_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_805_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_805_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_addr_0
    process(ptr_deref_105_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_base_resize
    process(arrayidx_103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_103;
      ov := iv(6 downto 0);
      ptr_deref_105_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_gather_scatter
    process(conv5212_80) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv5212_80;
      ov(15 downto 0) := iv;
      ptr_deref_105_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_root_address_inst
    process(ptr_deref_105_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_addr_0
    process(ptr_deref_122_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_base_resize
    process(iNsTr_13_119) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_119;
      ov := iv(6 downto 0);
      ptr_deref_122_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_gather_scatter
    process(ptr_deref_122_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_data_0;
      ov(15 downto 0) := iv;
      tmp1_123 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_root_address_inst
    process(ptr_deref_122_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_addr_0
    process(ptr_deref_171_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_171_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_171_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_base_resize
    process(iNsTr_5_169) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_169;
      ov := iv(6 downto 0);
      ptr_deref_171_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_gather_scatter
    process(conv5x_xlcssa_157) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv5x_xlcssa_157;
      ov(15 downto 0) := iv;
      ptr_deref_171_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_root_address_inst
    process(ptr_deref_171_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_171_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_171_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_addr_0
    process(ptr_deref_222_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_222_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_222_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_base_resize
    process(arrayidx21_213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx21_213;
      ov := iv(6 downto 0);
      ptr_deref_222_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_gather_scatter
    process(conv18_220) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv18_220;
      ov(15 downto 0) := iv;
      ptr_deref_222_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_root_address_inst
    process(ptr_deref_222_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_222_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_222_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_addr_0
    process(ptr_deref_239_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_239_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_base_resize
    process(iNsTr_21_236) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_236;
      ov := iv(6 downto 0);
      ptr_deref_239_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_gather_scatter
    process(ptr_deref_239_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_data_0;
      ov(15 downto 0) := iv;
      tmp12_240 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_root_address_inst
    process(ptr_deref_239_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_239_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_addr_0
    process(ptr_deref_290_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_290_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_290_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_base_resize
    process(arrayidx35_288) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35_288;
      ov := iv(0 downto 0);
      ptr_deref_290_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_gather_scatter
    process(conv32199_277) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv32199_277;
      ov(15 downto 0) := iv;
      ptr_deref_290_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_root_address_inst
    process(ptr_deref_290_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_290_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_290_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_addr_0
    process(ptr_deref_343_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_343_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_base_resize
    process(iNsTr_26_341) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_341;
      ov := iv(6 downto 0);
      ptr_deref_343_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_gather_scatter
    process(conv43_333) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_333;
      ov(15 downto 0) := iv;
      ptr_deref_343_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_root_address_inst
    process(ptr_deref_343_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_343_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_addr_0
    process(ptr_deref_362_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_362_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_362_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_base_resize
    process(iNsTr_29_360) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_360;
      ov := iv(6 downto 0);
      ptr_deref_362_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_gather_scatter
    process(conv45_352) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_352;
      ov(15 downto 0) := iv;
      ptr_deref_362_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_root_address_inst
    process(ptr_deref_362_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_362_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_362_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_addr_0
    process(ptr_deref_381_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_base_resize
    process(iNsTr_32_379) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_379;
      ov := iv(6 downto 0);
      ptr_deref_381_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_gather_scatter
    process(conv47_371) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv47_371;
      ov(15 downto 0) := iv;
      ptr_deref_381_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_root_address_inst
    process(ptr_deref_381_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_addr_0
    process(ptr_deref_394_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_base_resize
    process(iNsTr_34_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_391;
      ov := iv(6 downto 0);
      ptr_deref_394_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_gather_scatter
    process(ptr_deref_394_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_data_0;
      ov(15 downto 0) := iv;
      tmp49_395 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_root_address_inst
    process(ptr_deref_394_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_addr_0
    process(ptr_deref_410_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_410_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_base_resize
    process(iNsTr_35_407) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_407;
      ov := iv(6 downto 0);
      ptr_deref_410_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_gather_scatter
    process(ptr_deref_410_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_data_0;
      ov(15 downto 0) := iv;
      tmp51_411 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_root_address_inst
    process(ptr_deref_410_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_410_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_addr_0
    process(ptr_deref_426_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_base_resize
    process(iNsTr_36_423) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_423;
      ov := iv(6 downto 0);
      ptr_deref_426_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_gather_scatter
    process(ptr_deref_426_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_data_0;
      ov(15 downto 0) := iv;
      tmp53_427 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_root_address_inst
    process(ptr_deref_426_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_452_addr_0
    process(ptr_deref_452_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_452_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_452_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_452_base_resize
    process(iNsTr_37_449) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_449;
      ov := iv(6 downto 0);
      ptr_deref_452_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_452_gather_scatter
    process(ptr_deref_452_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_452_data_0;
      ov(15 downto 0) := iv;
      tmp57_453 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_452_root_address_inst
    process(ptr_deref_452_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_452_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_452_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_addr_0
    process(ptr_deref_468_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_base_resize
    process(iNsTr_38_465) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_465;
      ov := iv(6 downto 0);
      ptr_deref_468_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_gather_scatter
    process(ptr_deref_468_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_data_0;
      ov(15 downto 0) := iv;
      tmp59_469 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_root_address_inst
    process(ptr_deref_468_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_addr_0
    process(ptr_deref_47_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_base_resize
    process(iNsTr_1_45) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_45;
      ov := iv(6 downto 0);
      ptr_deref_47_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_gather_scatter
    process(conv_39) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_39;
      ov(15 downto 0) := iv;
      ptr_deref_47_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_root_address_inst
    process(ptr_deref_47_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_addr_0
    process(ptr_deref_484_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_484_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_base_resize
    process(iNsTr_39_481) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_481;
      ov := iv(6 downto 0);
      ptr_deref_484_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_gather_scatter
    process(ptr_deref_484_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_data_0;
      ov(15 downto 0) := iv;
      tmp62_485 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_root_address_inst
    process(ptr_deref_484_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_484_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_addr_0
    process(ptr_deref_500_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_500_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_base_resize
    process(iNsTr_40_497) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_497;
      ov := iv(6 downto 0);
      ptr_deref_500_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_gather_scatter
    process(ptr_deref_500_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_data_0;
      ov(15 downto 0) := iv;
      tmp65_501 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_root_address_inst
    process(ptr_deref_500_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_500_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_735_addr_0
    process(ptr_deref_735_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_735_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_735_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_735_base_resize
    process(arrayidx120_600) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx120_600;
      ov := iv(13 downto 0);
      ptr_deref_735_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_735_gather_scatter
    process(add116_733) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add116_733;
      ov(63 downto 0) := iv;
      ptr_deref_735_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_735_root_address_inst
    process(ptr_deref_735_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_735_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_735_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_addr_0
    process(ptr_deref_942_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_942_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_base_resize
    process(arrayidx181_807) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx181_807;
      ov := iv(10 downto 0);
      ptr_deref_942_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_gather_scatter
    process(add177_940) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add177_940;
      ov(63 downto 0) := iv;
      ptr_deref_942_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_root_address_inst
    process(ptr_deref_942_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_942_root_address <= ov(10 downto 0);
      --
    end process;
    if_stmt_143_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_135;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_143_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_143_branch_req_0,
          ack0 => if_stmt_143_branch_ack_0,
          ack1 => if_stmt_143_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_180_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp14203_179;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_180_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_180_branch_req_0,
          ack0 => if_stmt_180_branch_ack_0,
          ack1 => if_stmt_180_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_252_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp14_251;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_252_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_252_branch_req_0,
          ack0 => if_stmt_252_branch_ack_0,
          ack1 => if_stmt_252_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_312_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond6_311;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_312_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_312_branch_req_0,
          ack0 => if_stmt_312_branch_ack_0,
          ack1 => if_stmt_312_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_527_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp71192_526;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_527_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_527_branch_req_0,
          ack0 => if_stmt_527_branch_ack_0,
          ack1 => if_stmt_527_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_542_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp129189_541;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_542_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_542_branch_req_0,
          ack0 => if_stmt_542_branch_ack_0,
          ack1 => if_stmt_542_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_64_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp208_56;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_64_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_64_branch_req_0,
          ack0 => if_stmt_64_branch_ack_0,
          ack1 => if_stmt_64_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_749_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_748;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_749_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_749_branch_req_0,
          ack0 => if_stmt_749_branch_ack_0,
          ack1 => if_stmt_749_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_955;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_956_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_956_branch_req_0,
          ack0 => if_stmt_956_branch_ack_0,
          ack1 => if_stmt_956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_565_inst
    process(tmp233_554) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp233_554, type_cast_564_wire_constant, tmp_var);
      tmp233x_xop_566 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_772_inst
    process(tmp221_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp221_761, type_cast_771_wire_constant, tmp_var);
      tmp221x_xop_773 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_112_inst
    process(indvar249_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar249_73, type_cast_111_wire_constant, tmp_var);
      tmp251_113 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_201_inst
    process(indvar244_189) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar244_189, type_cast_200_wire_constant, tmp_var);
      tmp3_202 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_229_inst
    process(indvar244_189) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar244_189, type_cast_228_wire_constant, tmp_var);
      tmp246_230 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_304_inst
    process(indvar241_270) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar241_270, type_cast_303_wire_constant, tmp_var);
      indvarx_xnext242_305 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_575_inst
    process(iNsTr_43_570) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_43_570, type_cast_574_wire_constant, tmp_var);
      xx_xop253_576 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_742_inst
    process(indvar226_586) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar226_586, type_cast_741_wire_constant, tmp_var);
      indvarx_xnext227_743 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_782_inst
    process(iNsTr_56_777) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_56_777, type_cast_781_wire_constant, tmp_var);
      xx_xop_783 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_91_inst
    process(indvar249_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar249_73, type_cast_90_wire_constant, tmp_var);
      tmp_92 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_949_inst
    process(indvar_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_793, type_cast_948_wire_constant, tmp_var);
      indvarx_xnext_950 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_178_inst
    process(conv5x_xlcssa_157) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv5x_xlcssa_157, type_cast_177_wire_constant, tmp_var);
      cmp14203_179 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_310_inst
    process(indvarx_xnext242_305) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext242_305, type_cast_309_wire_constant, tmp_var);
      exitcond6_311 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_747_inst
    process(indvarx_xnext227_743, tmp238_583) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext227_743, tmp238_583, tmp_var);
      exitcond_748 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_954_inst
    process(indvarx_xnext_950, tmp225_790) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_950, tmp225_790, tmp_var);
      exitcond5_955 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_54_inst
    process(call_35) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_35, type_cast_53_wire_constant, tmp_var);
      cmp208_56 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_553_inst
    process(mul55_441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul55_441, type_cast_552_wire_constant, tmp_var);
      tmp233_554 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_760_inst
    process(mul67_520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul67_520, type_cast_759_wire_constant, tmp_var);
      tmp221_761 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_435_inst
    process(conv52_415, conv50_399) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv52_415, conv50_399, tmp_var);
      mul_436 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_440_inst
    process(mul_436, conv54_431) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_436, conv54_431, tmp_var);
      mul55_441 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_509_inst
    process(conv60_473, conv58_457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv60_473, conv58_457, tmp_var);
      mul61_510 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_514_inst
    process(mul61_510, conv63_489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul61_510, conv63_489, tmp_var);
      mul64_515 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_519_inst
    process(mul64_515, conv66_505) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul64_515, conv66_505, tmp_var);
      mul67_520 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_624_inst
    process(shl_613, conv80_620) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_613, conv80_620, tmp_var);
      add_625 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_642_inst
    process(shl82_631, conv85_638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl82_631, conv85_638, tmp_var);
      add86_643 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_660_inst
    process(shl88_649, conv91_656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_649, conv91_656, tmp_var);
      add92_661 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_678_inst
    process(shl94_667, conv97_674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_667, conv97_674, tmp_var);
      add98_679 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_696_inst
    process(shl100_685, conv103_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_685, conv103_692, tmp_var);
      add104_697 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_714_inst
    process(shl106_703, conv109_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_703, conv109_710, tmp_var);
      add110_715 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_732_inst
    process(shl112_721, conv115_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl112_721, conv115_728, tmp_var);
      add116_733 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_831_inst
    process(shl137_820, conv140_827) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl137_820, conv140_827, tmp_var);
      add141_832 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_849_inst
    process(shl143_838, conv146_845) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl143_838, conv146_845, tmp_var);
      add147_850 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_867_inst
    process(shl149_856, conv152_863) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl149_856, conv152_863, tmp_var);
      add153_868 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_885_inst
    process(shl155_874, conv158_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl155_874, conv158_881, tmp_var);
      add159_886 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_903_inst
    process(shl161_892, conv164_899) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl161_892, conv164_899, tmp_var);
      add165_904 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_921_inst
    process(shl167_910, conv170_917) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_910, conv170_917, tmp_var);
      add171_922 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_939_inst
    process(shl173_928, conv176_935) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_928, conv176_935, tmp_var);
      add177_940 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_612_inst
    process(conv76_607) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv76_607, type_cast_611_wire_constant, tmp_var);
      shl_613 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_630_inst
    process(add_625) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_625, type_cast_629_wire_constant, tmp_var);
      shl82_631 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_648_inst
    process(add86_643) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add86_643, type_cast_647_wire_constant, tmp_var);
      shl88_649 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_666_inst
    process(add92_661) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_661, type_cast_665_wire_constant, tmp_var);
      shl94_667 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_684_inst
    process(add98_679) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_679, type_cast_683_wire_constant, tmp_var);
      shl100_685 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_702_inst
    process(add104_697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_697, type_cast_701_wire_constant, tmp_var);
      shl106_703 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_720_inst
    process(add110_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add110_715, type_cast_719_wire_constant, tmp_var);
      shl112_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_819_inst
    process(conv135_814) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv135_814, type_cast_818_wire_constant, tmp_var);
      shl137_820 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_837_inst
    process(add141_832) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add141_832, type_cast_836_wire_constant, tmp_var);
      shl143_838 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_855_inst
    process(add147_850) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add147_850, type_cast_854_wire_constant, tmp_var);
      shl149_856 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_873_inst
    process(add153_868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add153_868, type_cast_872_wire_constant, tmp_var);
      shl155_874 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_891_inst
    process(add159_886) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add159_886, type_cast_890_wire_constant, tmp_var);
      shl161_892 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_909_inst
    process(add165_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add165_904, type_cast_908_wire_constant, tmp_var);
      shl167_910 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_927_inst
    process(add171_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_922, type_cast_926_wire_constant, tmp_var);
      shl173_928 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_134_inst
    process(type_cast_131_wire, type_cast_133_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_131_wire, type_cast_133_wire, tmp_var);
      cmp_135 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_250_inst
    process(type_cast_247_wire, type_cast_249_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_247_wire, type_cast_249_wire, tmp_var);
      cmp14_251 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_525_inst
    process(mul55_441) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul55_441, type_cast_524_wire_constant, tmp_var);
      cmp71192_526 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_540_inst
    process(mul67_520) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul67_520, type_cast_539_wire_constant, tmp_var);
      cmp129189_541 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_559_inst
    process(tmp233_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp233_554, type_cast_558_wire_constant, tmp_var);
      tmp234_560 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_766_inst
    process(tmp221_761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp221_761, type_cast_765_wire_constant, tmp_var);
      tmp222_767 <= tmp_var; --
    end process;
    -- shared split operator group (57) : array_obj_ref_101_index_offset 
    ApIntAdd_group_57: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar249_100_scaled;
      array_obj_ref_101_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_101_index_offset_req_0;
      array_obj_ref_101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_101_index_offset_req_1;
      array_obj_ref_101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_57_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : array_obj_ref_211_index_offset 
    ApIntAdd_group_58: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar244_210_scaled;
      array_obj_ref_211_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_211_index_offset_req_0;
      array_obj_ref_211_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_211_index_offset_req_1;
      array_obj_ref_211_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_58_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : array_obj_ref_598_index_offset 
    ApIntAdd_group_59: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar226_597_scaled;
      array_obj_ref_598_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_598_index_offset_req_0;
      array_obj_ref_598_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_598_index_offset_req_1;
      array_obj_ref_598_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_59_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_59_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : array_obj_ref_805_index_offset 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_804_scaled;
      array_obj_ref_805_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_805_index_offset_req_0;
      array_obj_ref_805_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_805_index_offset_req_1;
      array_obj_ref_805_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared load operator group (0) : ptr_deref_122_load_0 ptr_deref_394_load_0 ptr_deref_410_load_0 ptr_deref_426_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_122_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_394_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_410_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_426_load_0_req_0;
      ptr_deref_122_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_394_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_410_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_426_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_122_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_394_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_410_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_426_load_0_req_1;
      ptr_deref_122_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_394_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_410_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_426_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_122_word_address_0 & ptr_deref_394_word_address_0 & ptr_deref_410_word_address_0 & ptr_deref_426_word_address_0;
      ptr_deref_122_data_0 <= data_out(63 downto 48);
      ptr_deref_394_data_0 <= data_out(47 downto 32);
      ptr_deref_410_data_0 <= data_out(31 downto 16);
      ptr_deref_426_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_239_load_0 ptr_deref_452_load_0 ptr_deref_468_load_0 ptr_deref_484_load_0 ptr_deref_500_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_239_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_452_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_468_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_484_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_500_load_0_req_0;
      ptr_deref_239_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_452_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_468_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_484_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_500_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_239_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_452_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_468_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_484_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_500_load_0_req_1;
      ptr_deref_239_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_452_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_468_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_484_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_500_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_239_word_address_0 & ptr_deref_452_word_address_0 & ptr_deref_468_word_address_0 & ptr_deref_484_word_address_0 & ptr_deref_500_word_address_0;
      ptr_deref_239_data_0 <= data_out(79 downto 64);
      ptr_deref_452_data_0 <= data_out(63 downto 48);
      ptr_deref_468_data_0 <= data_out(47 downto 32);
      ptr_deref_484_data_0 <= data_out(31 downto 16);
      ptr_deref_500_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : STORE_padding_324_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_324_store_0_req_0;
      STORE_padding_324_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_324_store_0_req_1;
      STORE_padding_324_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_324_word_address_0;
      data_in <= STORE_padding_324_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_47_store_0 ptr_deref_105_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_47_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_105_store_0_req_0;
      ptr_deref_47_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_105_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_47_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_105_store_0_req_1;
      ptr_deref_47_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_105_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_47_word_address_0 & ptr_deref_105_word_address_0;
      data_in <= ptr_deref_47_data_0 & ptr_deref_105_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(15 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_222_store_0 ptr_deref_171_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_222_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_171_store_0_req_0;
      ptr_deref_222_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_171_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_222_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_171_store_0_req_1;
      ptr_deref_222_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_171_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_222_word_address_0 & ptr_deref_171_word_address_0;
      data_in <= ptr_deref_222_data_0 & ptr_deref_171_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(15 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_290_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_290_store_0_req_0;
      ptr_deref_290_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_290_store_0_req_1;
      ptr_deref_290_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_290_word_address_0;
      data_in <= ptr_deref_290_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_343_store_0 ptr_deref_362_store_0 ptr_deref_381_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_343_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_362_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_381_store_0_req_0;
      ptr_deref_343_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_362_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_381_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_343_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_362_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_381_store_0_req_1;
      ptr_deref_343_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_362_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_381_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_343_word_address_0 & ptr_deref_362_word_address_0 & ptr_deref_381_word_address_0;
      data_in <= ptr_deref_343_data_0 & ptr_deref_362_data_0 & ptr_deref_381_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(15 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_735_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_735_store_0_req_0;
      ptr_deref_735_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_735_store_0_req_1;
      ptr_deref_735_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_735_word_address_0;
      data_in <= ptr_deref_735_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_942_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_942_store_0_req_0;
      ptr_deref_942_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_942_store_0_req_1;
      ptr_deref_942_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_942_word_address_0;
      data_in <= ptr_deref_942_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(10 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_651_inst RPIPE_ConvTranspose_input_pipe_615_inst RPIPE_ConvTranspose_input_pipe_602_inst RPIPE_ConvTranspose_input_pipe_633_inst RPIPE_ConvTranspose_input_pipe_262_inst RPIPE_ConvTranspose_input_pipe_294_inst RPIPE_ConvTranspose_input_pipe_137_inst RPIPE_ConvTranspose_input_pipe_215_inst RPIPE_ConvTranspose_input_pipe_876_inst RPIPE_ConvTranspose_input_pipe_669_inst RPIPE_ConvTranspose_input_pipe_687_inst RPIPE_ConvTranspose_input_pipe_705_inst RPIPE_ConvTranspose_input_pipe_894_inst RPIPE_ConvTranspose_input_pipe_723_inst RPIPE_ConvTranspose_input_pipe_912_inst RPIPE_ConvTranspose_input_pipe_930_inst RPIPE_ConvTranspose_input_pipe_809_inst RPIPE_ConvTranspose_input_pipe_822_inst RPIPE_ConvTranspose_input_pipe_840_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_58_inst RPIPE_ConvTranspose_input_pipe_328_inst RPIPE_ConvTranspose_input_pipe_347_inst RPIPE_ConvTranspose_input_pipe_366_inst RPIPE_ConvTranspose_input_pipe_858_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_651_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_615_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_602_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_633_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_137_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_215_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_669_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_687_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_930_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_809_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_822_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_840_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_651_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_615_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_602_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_633_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_137_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_215_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_669_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_687_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_930_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_809_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_822_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_840_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_651_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_615_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_602_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_633_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_137_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_215_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_876_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_669_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_687_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_894_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_912_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_930_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_809_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_822_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_840_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_858_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_651_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_615_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_602_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_633_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_137_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_215_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_876_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_669_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_687_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_894_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_912_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_930_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_809_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_822_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_840_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_858_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call89_652 <= data_out(199 downto 192);
      call78_616 <= data_out(191 downto 184);
      call75_603 <= data_out(183 downto 176);
      call83_634 <= data_out(175 downto 168);
      call31196_263 <= data_out(167 downto 160);
      call31_295 <= data_out(159 downto 152);
      call4_138 <= data_out(151 downto 144);
      call17_216 <= data_out(143 downto 136);
      call156_877 <= data_out(135 downto 128);
      call95_670 <= data_out(127 downto 120);
      call101_688 <= data_out(119 downto 112);
      call107_706 <= data_out(111 downto 104);
      call162_895 <= data_out(103 downto 96);
      call113_724 <= data_out(95 downto 88);
      call168_913 <= data_out(87 downto 80);
      call174_931 <= data_out(79 downto 72);
      call134_810 <= data_out(71 downto 64);
      call138_823 <= data_out(63 downto 56);
      call144_841 <= data_out(55 downto 48);
      call_35 <= data_out(47 downto 40);
      call4209_59 <= data_out(39 downto 32);
      call42_329 <= data_out(31 downto 24);
      call44_348 <= data_out(23 downto 16);
      call46_367 <= data_out(15 downto 8);
      call150_859 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(99 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(55 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(75 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 21),
      memory_space_0_lr_tag => memory_space_0_lr_tag(83 downto 63),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 48),
      memory_space_0_lc_tag => memory_space_0_lc_tag(11 downto 9),
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 48),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(79 downto 60),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 48),
      memory_space_2_lc_tag => memory_space_2_lc_tag(7 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(55 downto 42),
      memory_space_3_lr_tag => memory_space_3_lr_tag(75 downto 57),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(255 downto 192),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 3),
      memory_space_6_lr_req => memory_space_6_lr_req(3 downto 3),
      memory_space_6_lr_ack => memory_space_6_lr_ack(3 downto 3),
      memory_space_6_lr_addr => memory_space_6_lr_addr(3 downto 3),
      memory_space_6_lr_tag => memory_space_6_lr_tag(75 downto 57),
      memory_space_6_lc_req => memory_space_6_lc_req(3 downto 3),
      memory_space_6_lc_ack => memory_space_6_lc_ack(3 downto 3),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 48),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(79 downto 60),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 6),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(55 downto 42),
      memory_space_5_sr_data => memory_space_5_sr_data(255 downto 192),
      memory_space_5_sr_tag => memory_space_5_sr_tag(75 downto 57),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(20 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(62 downto 42),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(47 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(8 downto 6),
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(47 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(59 downto 40),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(47 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 4),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(56 downto 38),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 2),
      memory_space_6_lr_req => memory_space_6_lr_req(2 downto 2),
      memory_space_6_lr_ack => memory_space_6_lr_ack(2 downto 2),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 2),
      memory_space_6_lr_tag => memory_space_6_lr_tag(56 downto 38),
      memory_space_6_lc_req => memory_space_6_lc_req(2 downto 2),
      memory_space_6_lc_ack => memory_space_6_lc_ack(2 downto 2),
      memory_space_6_lc_data => memory_space_6_lc_data(47 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(59 downto 40),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(5 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(41 downto 28),
      memory_space_5_sr_data => memory_space_5_sr_data(191 downto 128),
      memory_space_5_sr_tag => memory_space_5_sr_tag(56 downto 38),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 7),
      memory_space_0_lr_tag => memory_space_0_lr_tag(41 downto 21),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 16),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 16),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(39 downto 20),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 16),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 1),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(37 downto 19),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 16),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(39 downto 20),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 2),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(27 downto 14),
      memory_space_5_sr_data => memory_space_5_sr_data(127 downto 64),
      memory_space_5_sr_tag => memory_space_5_sr_tag(37 downto 19),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(15 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(15 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(19 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(13 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(99 downto 80),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(79 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 8),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(4 downto 4),
      memory_space_0_lr_ack => memory_space_0_lr_ack(4 downto 4),
      memory_space_0_lr_addr => memory_space_0_lr_addr(34 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(104 downto 84),
      memory_space_0_lc_req => memory_space_0_lc_req(4 downto 4),
      memory_space_0_lc_ack => memory_space_0_lc_ack(4 downto 4),
      memory_space_0_lc_data => memory_space_0_lc_data(79 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(14 downto 12),
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(79 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(15 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(10 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(0 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(19 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 4,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
